library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package PkgLUT is
  -- Layer 0 
  subtype  lut_array_t_0 is array (0 to 63) of signed(4 downto 0);

  constant LUT_0_0_0_DATA : lut_array_t_0 := (
    0 => "00010", --    2
    1 => "00011", --    3
    2 => "00011", --    3
    3 => "00011", --    3
    4 => "00011", --    3
    5 => "00011", --    3
    6 => "00011", --    3
    7 => "00011", --    3
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11110", --   -2
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00100", --    4
    63 => "00100", --    4
  );

  constant LUT_0_0_1_DATA : lut_array_t_0 := (
    0 => "00011", --    3
    1 => "00011", --    3
    2 => "00011", --    3
    3 => "00011", --    3
    4 => "00011", --    3
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00001", --    1
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "11111", --   -1
    11 => "11110", --   -2
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11100", --   -4
    15 => "11100", --   -4
    16 => "11100", --   -4
    17 => "11100", --   -4
    18 => "11100", --   -4
    19 => "11100", --   -4
    20 => "11100", --   -4
    21 => "11100", --   -4
    22 => "11100", --   -4
    23 => "11101", --   -3
    24 => "11101", --   -3
    25 => "11101", --   -3
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11111", --   -1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00010", --    2
    36 => "00011", --    3
    37 => "00011", --    3
    38 => "00011", --    3
    39 => "00100", --    4
    40 => "00100", --    4
    41 => "00100", --    4
    42 => "00101", --    5
    43 => "00101", --    5
    44 => "00101", --    5
    45 => "00110", --    6
    46 => "00110", --    6
    47 => "00110", --    6
    48 => "00111", --    7
    49 => "00111", --    7
    50 => "01000", --    8
    51 => "01000", --    8
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01010", --   10
    57 => "01011", --   11
    58 => "01011", --   11
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01100", --   12
    62 => "01101", --   13
    63 => "01101", --   13
  );

  constant LUT_0_0_2_DATA : lut_array_t_0 := (
    0 => "00101", --    5
    1 => "00110", --    6
    2 => "00110", --    6
    3 => "00110", --    6
    4 => "00110", --    6
    5 => "00101", --    5
    6 => "00101", --    5
    7 => "00101", --    5
    8 => "00100", --    4
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00100", --    4
    20 => "00100", --    4
    21 => "00100", --    4
    22 => "00100", --    4
    23 => "00011", --    3
    24 => "00011", --    3
    25 => "00011", --    3
    26 => "00011", --    3
    27 => "00010", --    2
    28 => "00010", --    2
    29 => "00010", --    2
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11110", --   -2
    37 => "11101", --   -3
    38 => "11101", --   -3
    39 => "11100", --   -4
    40 => "11100", --   -4
    41 => "11011", --   -5
    42 => "11010", --   -6
    43 => "11001", --   -7
    44 => "11001", --   -7
    45 => "11000", --   -8
    46 => "10111", --   -9
    47 => "10110", --  -10
    48 => "10110", --  -10
    49 => "10101", --  -11
    50 => "10100", --  -12
    51 => "10100", --  -12
    52 => "10011", --  -13
    53 => "10010", --  -14
    54 => "10010", --  -14
    55 => "10001", --  -15
    56 => "10001", --  -15
    57 => "10000", --  -16
    58 => "10000", --  -16
    59 => "10000", --  -16
    60 => "10000", --  -16
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_0_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00010", --    2
    25 => "00010", --    2
    26 => "00010", --    2
    27 => "00010", --    2
    28 => "00010", --    2
    29 => "00010", --    2
    30 => "00010", --    2
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11101", --   -3
    44 => "11101", --   -3
    45 => "11100", --   -4
    46 => "11100", --   -4
    47 => "11011", --   -5
    48 => "11011", --   -5
    49 => "11010", --   -6
    50 => "11010", --   -6
    51 => "11001", --   -7
    52 => "11001", --   -7
    53 => "11000", --   -8
    54 => "11000", --   -8
    55 => "11000", --   -8
    56 => "10111", --   -9
    57 => "10111", --   -9
    58 => "10111", --   -9
    59 => "10111", --   -9
    60 => "10111", --   -9
    61 => "10111", --   -9
    62 => "10110", --  -10
    63 => "10110", --  -10
  );

  constant LUT_0_0_4_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11101", --   -3
    3 => "11101", --   -3
    4 => "11101", --   -3
    5 => "11100", --   -4
    6 => "11100", --   -4
    7 => "11011", --   -5
    8 => "11011", --   -5
    9 => "11010", --   -6
    10 => "11010", --   -6
    11 => "11001", --   -7
    12 => "11001", --   -7
    13 => "11001", --   -7
    14 => "11001", --   -7
    15 => "11000", --   -8
    16 => "11000", --   -8
    17 => "11001", --   -7
    18 => "11001", --   -7
    19 => "11001", --   -7
    20 => "11001", --   -7
    21 => "11010", --   -6
    22 => "11010", --   -6
    23 => "11010", --   -6
    24 => "11011", --   -5
    25 => "11100", --   -4
    26 => "11100", --   -4
    27 => "11101", --   -3
    28 => "11110", --   -2
    29 => "11110", --   -2
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00001", --    1
    34 => "00010", --    2
    35 => "00011", --    3
    36 => "00011", --    3
    37 => "00100", --    4
    38 => "00101", --    5
    39 => "00110", --    6
    40 => "00110", --    6
    41 => "00111", --    7
    42 => "01000", --    8
    43 => "01001", --    9
    44 => "01010", --   10
    45 => "01010", --   10
    46 => "01011", --   11
    47 => "01100", --   12
    48 => "01100", --   12
    49 => "01101", --   13
    50 => "01101", --   13
    51 => "01110", --   14
    52 => "01110", --   14
    53 => "01111", --   15
    54 => "01111", --   15
    55 => "01111", --   15
    56 => "01111", --   15
    57 => "01111", --   15
    58 => "01111", --   15
    59 => "01111", --   15
    60 => "01111", --   15
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_0_5_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00001", --    1
    60 => "00001", --    1
    61 => "00001", --    1
    62 => "00001", --    1
    63 => "00001", --    1
  );

  constant LUT_0_0_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "00000", --    0
    58 => "00000", --    0
    59 => "00000", --    0
    60 => "00000", --    0
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_0_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11101", --   -3
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11100", --   -4
    53 => "11100", --   -4
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11100", --   -4
    57 => "11100", --   -4
    58 => "11011", --   -5
    59 => "11011", --   -5
    60 => "11011", --   -5
    61 => "11011", --   -5
    62 => "11010", --   -6
    63 => "11010", --   -6
  );

  constant LUT_0_1_0_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00100", --    4
    47 => "00101", --    5
    48 => "00101", --    5
    49 => "00101", --    5
    50 => "00110", --    6
    51 => "00110", --    6
    52 => "00110", --    6
    53 => "00110", --    6
    54 => "00111", --    7
    55 => "00111", --    7
    56 => "00111", --    7
    57 => "01000", --    8
    58 => "01000", --    8
    59 => "01000", --    8
    60 => "01000", --    8
    61 => "01001", --    9
    62 => "01001", --    9
    63 => "01010", --   10
  );

  constant LUT_0_1_1_DATA : lut_array_t_0 := (
    0 => "11011", --   -5
    1 => "11011", --   -5
    2 => "11011", --   -5
    3 => "11011", --   -5
    4 => "11011", --   -5
    5 => "11100", --   -4
    6 => "11100", --   -4
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11101", --   -3
    19 => "11101", --   -3
    20 => "11101", --   -3
    21 => "11101", --   -3
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00011", --    3
    39 => "00011", --    3
    40 => "00100", --    4
    41 => "00101", --    5
    42 => "00101", --    5
    43 => "00110", --    6
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "01000", --    8
    47 => "01000", --    8
    48 => "01001", --    9
    49 => "01001", --    9
    50 => "01001", --    9
    51 => "01010", --   10
    52 => "01010", --   10
    53 => "01010", --   10
    54 => "01011", --   11
    55 => "01011", --   11
    56 => "01011", --   11
    57 => "01100", --   12
    58 => "01100", --   12
    59 => "01101", --   13
    60 => "01101", --   13
    61 => "01110", --   14
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_1_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11101", --   -3
    58 => "11101", --   -3
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_1_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "00000", --    0
    58 => "00000", --    0
    59 => "00000", --    0
    60 => "00000", --    0
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_1_4_DATA : lut_array_t_0 := (
    0 => "11011", --   -5
    1 => "11011", --   -5
    2 => "11011", --   -5
    3 => "11011", --   -5
    4 => "11011", --   -5
    5 => "11011", --   -5
    6 => "11100", --   -4
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11110", --   -2
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00010", --    2
    35 => "00010", --    2
    36 => "00011", --    3
    37 => "00011", --    3
    38 => "00011", --    3
    39 => "00011", --    3
    40 => "00100", --    4
    41 => "00100", --    4
    42 => "00100", --    4
    43 => "00100", --    4
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00100", --    4
    47 => "00100", --    4
    48 => "00100", --    4
    49 => "00100", --    4
    50 => "00100", --    4
    51 => "00100", --    4
    52 => "00100", --    4
    53 => "00100", --    4
    54 => "00101", --    5
    55 => "00101", --    5
    56 => "00110", --    6
    57 => "00110", --    6
    58 => "00111", --    7
    59 => "00111", --    7
    60 => "01000", --    8
    61 => "01000", --    8
    62 => "01001", --    9
    63 => "01001", --    9
  );

  constant LUT_0_1_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00101", --    5
    47 => "00101", --    5
    48 => "00110", --    6
    49 => "00110", --    6
    50 => "00111", --    7
    51 => "00111", --    7
    52 => "00111", --    7
    53 => "00111", --    7
    54 => "01000", --    8
    55 => "01000", --    8
    56 => "01000", --    8
    57 => "01000", --    8
    58 => "01000", --    8
    59 => "01000", --    8
    60 => "01000", --    8
    61 => "01001", --    9
    62 => "01001", --    9
    63 => "01001", --    9
  );

  constant LUT_0_1_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "00000", --    0
    58 => "00000", --    0
    59 => "00000", --    0
    60 => "00000", --    0
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_1_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00100", --    4
    53 => "00100", --    4
    54 => "00100", --    4
    55 => "00100", --    4
    56 => "00101", --    5
    57 => "00101", --    5
    58 => "00101", --    5
    59 => "00101", --    5
    60 => "00101", --    5
    61 => "00110", --    6
    62 => "00110", --    6
    63 => "00110", --    6
  );

  constant LUT_0_2_0_DATA : lut_array_t_0 := (
    0 => "00010", --    2
    1 => "00010", --    2
    2 => "00011", --    3
    3 => "00011", --    3
    4 => "00011", --    3
    5 => "00011", --    3
    6 => "00100", --    4
    7 => "00100", --    4
    8 => "00100", --    4
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00101", --    5
    12 => "00101", --    5
    13 => "00101", --    5
    14 => "00100", --    4
    15 => "00100", --    4
    16 => "00100", --    4
    17 => "00100", --    4
    18 => "00011", --    3
    19 => "00011", --    3
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00000", --    0
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11110", --   -2
    31 => "11110", --   -2
    32 => "11110", --   -2
    33 => "11110", --   -2
    34 => "11110", --   -2
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11101", --   -3
    43 => "11101", --   -3
    44 => "11100", --   -4
    45 => "11100", --   -4
    46 => "11100", --   -4
    47 => "11100", --   -4
    48 => "11011", --   -5
    49 => "11011", --   -5
    50 => "11011", --   -5
    51 => "11010", --   -6
    52 => "11010", --   -6
    53 => "11001", --   -7
    54 => "11001", --   -7
    55 => "11000", --   -8
    56 => "11000", --   -8
    57 => "10111", --   -9
    58 => "10111", --   -9
    59 => "10110", --  -10
    60 => "10110", --  -10
    61 => "10110", --  -10
    62 => "10110", --  -10
    63 => "10110", --  -10
  );

  constant LUT_0_2_1_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00011", --    3
    9 => "00011", --    3
    10 => "00011", --    3
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00011", --    3
    20 => "00011", --    3
    21 => "00011", --    3
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00010", --    2
    25 => "00010", --    2
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11101", --   -3
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11100", --   -4
    43 => "11100", --   -4
    44 => "11011", --   -5
    45 => "11011", --   -5
    46 => "11010", --   -6
    47 => "11001", --   -7
    48 => "11001", --   -7
    49 => "11000", --   -8
    50 => "10111", --   -9
    51 => "10111", --   -9
    52 => "10110", --  -10
    53 => "10101", --  -11
    54 => "10100", --  -12
    55 => "10100", --  -12
    56 => "10011", --  -13
    57 => "10010", --  -14
    58 => "10010", --  -14
    59 => "10001", --  -15
    60 => "10001", --  -15
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_2_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00010", --    2
    25 => "00010", --    2
    26 => "00010", --    2
    27 => "00010", --    2
    28 => "00010", --    2
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11100", --   -4
    41 => "11100", --   -4
    42 => "11011", --   -5
    43 => "11011", --   -5
    44 => "11011", --   -5
    45 => "11011", --   -5
    46 => "11011", --   -5
    47 => "11010", --   -6
    48 => "11010", --   -6
    49 => "11010", --   -6
    50 => "11010", --   -6
    51 => "11010", --   -6
    52 => "11010", --   -6
    53 => "11010", --   -6
    54 => "11010", --   -6
    55 => "11001", --   -7
    56 => "11001", --   -7
    57 => "11001", --   -7
    58 => "11000", --   -8
    59 => "11000", --   -8
    60 => "10111", --   -9
    61 => "10111", --   -9
    62 => "10111", --   -9
    63 => "10110", --  -10
  );

  constant LUT_0_2_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00011", --    3
    46 => "00011", --    3
    47 => "00100", --    4
    48 => "00100", --    4
    49 => "00100", --    4
    50 => "00101", --    5
    51 => "00101", --    5
    52 => "00101", --    5
    53 => "00110", --    6
    54 => "00110", --    6
    55 => "00110", --    6
    56 => "00110", --    6
    57 => "00111", --    7
    58 => "00111", --    7
    59 => "00111", --    7
    60 => "00111", --    7
    61 => "00111", --    7
    62 => "00111", --    7
    63 => "00111", --    7
  );

  constant LUT_0_2_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00010", --    2
    63 => "00010", --    2
  );

  constant LUT_0_2_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00011", --    3
    41 => "00011", --    3
    42 => "00100", --    4
    43 => "00100", --    4
    44 => "00101", --    5
    45 => "00101", --    5
    46 => "00110", --    6
    47 => "00110", --    6
    48 => "00110", --    6
    49 => "00111", --    7
    50 => "00111", --    7
    51 => "01000", --    8
    52 => "01000", --    8
    53 => "01000", --    8
    54 => "01001", --    9
    55 => "01001", --    9
    56 => "01010", --   10
    57 => "01011", --   11
    58 => "01011", --   11
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01101", --   13
    62 => "01110", --   14
    63 => "01110", --   14
  );

  constant LUT_0_2_6_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11101", --   -3
    6 => "11101", --   -3
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11011", --   -5
    10 => "11010", --   -6
    11 => "11010", --   -6
    12 => "11010", --   -6
    13 => "11001", --   -7
    14 => "11001", --   -7
    15 => "11010", --   -6
    16 => "11010", --   -6
    17 => "11010", --   -6
    18 => "11010", --   -6
    19 => "11011", --   -5
    20 => "11011", --   -5
    21 => "11100", --   -4
    22 => "11100", --   -4
    23 => "11100", --   -4
    24 => "11101", --   -3
    25 => "11101", --   -3
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11110", --   -2
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00011", --    3
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00101", --    5
    47 => "00101", --    5
    48 => "00110", --    6
    49 => "00110", --    6
    50 => "00111", --    7
    51 => "01000", --    8
    52 => "01000", --    8
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01011", --   11
    57 => "01011", --   11
    58 => "01011", --   11
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01100", --   12
    62 => "01100", --   12
    63 => "01100", --   12
  );

  constant LUT_0_2_7_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11101", --   -3
    3 => "11101", --   -3
    4 => "11101", --   -3
    5 => "11101", --   -3
    6 => "11100", --   -4
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11100", --   -4
    12 => "11100", --   -4
    13 => "11100", --   -4
    14 => "11100", --   -4
    15 => "11100", --   -4
    16 => "11100", --   -4
    17 => "11100", --   -4
    18 => "11100", --   -4
    19 => "11100", --   -4
    20 => "11100", --   -4
    21 => "11101", --   -3
    22 => "11101", --   -3
    23 => "11101", --   -3
    24 => "11101", --   -3
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00010", --    2
    36 => "00010", --    2
    37 => "00011", --    3
    38 => "00011", --    3
    39 => "00100", --    4
    40 => "00100", --    4
    41 => "00101", --    5
    42 => "00101", --    5
    43 => "00110", --    6
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "01000", --    8
    47 => "01001", --    9
    48 => "01001", --    9
    49 => "01010", --   10
    50 => "01011", --   11
    51 => "01011", --   11
    52 => "01100", --   12
    53 => "01100", --   12
    54 => "01101", --   13
    55 => "01101", --   13
    56 => "01110", --   14
    57 => "01110", --   14
    58 => "01111", --   15
    59 => "01111", --   15
    60 => "01111", --   15
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_3_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11101", --   -3
    25 => "11101", --   -3
    26 => "11101", --   -3
    27 => "11101", --   -3
    28 => "11101", --   -3
    29 => "11110", --   -2
    30 => "11110", --   -2
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00011", --    3
    47 => "00011", --    3
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_3_1_DATA : lut_array_t_0 := (
    0 => "00010", --    2
    1 => "00011", --    3
    2 => "00011", --    3
    3 => "00011", --    3
    4 => "00100", --    4
    5 => "00100", --    4
    6 => "00100", --    4
    7 => "00101", --    5
    8 => "00101", --    5
    9 => "00101", --    5
    10 => "00110", --    6
    11 => "00110", --    6
    12 => "00110", --    6
    13 => "00110", --    6
    14 => "00110", --    6
    15 => "00111", --    7
    16 => "00111", --    7
    17 => "00111", --    7
    18 => "00111", --    7
    19 => "00111", --    7
    20 => "00111", --    7
    21 => "00111", --    7
    22 => "00111", --    7
    23 => "00110", --    6
    24 => "00110", --    6
    25 => "00101", --    5
    26 => "00101", --    5
    27 => "00100", --    4
    28 => "00010", --    2
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "11111", --   -1
    32 => "11110", --   -2
    33 => "11100", --   -4
    34 => "11011", --   -5
    35 => "11010", --   -6
    36 => "11001", --   -7
    37 => "11001", --   -7
    38 => "11000", --   -8
    39 => "10111", --   -9
    40 => "10111", --   -9
    41 => "10111", --   -9
    42 => "10111", --   -9
    43 => "10111", --   -9
    44 => "10111", --   -9
    45 => "10111", --   -9
    46 => "10111", --   -9
    47 => "10111", --   -9
    48 => "10111", --   -9
    49 => "10111", --   -9
    50 => "10111", --   -9
    51 => "10110", --  -10
    52 => "10110", --  -10
    53 => "10110", --  -10
    54 => "10101", --  -11
    55 => "10101", --  -11
    56 => "10100", --  -12
    57 => "10011", --  -13
    58 => "10011", --  -13
    59 => "10010", --  -14
    60 => "10001", --  -15
    61 => "10001", --  -15
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_3_2_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11101", --   -3
    57 => "11101", --   -3
    58 => "11101", --   -3
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_3_3_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11110", --   -2
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00010", --    2
    37 => "00011", --    3
    38 => "00011", --    3
    39 => "00100", --    4
    40 => "00101", --    5
    41 => "00101", --    5
    42 => "00110", --    6
    43 => "00111", --    7
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "01000", --    8
    47 => "01000", --    8
    48 => "01000", --    8
    49 => "01000", --    8
    50 => "01000", --    8
    51 => "01001", --    9
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01011", --   11
    57 => "01011", --   11
    58 => "01100", --   12
    59 => "01100", --   12
    60 => "01101", --   13
    61 => "01110", --   14
    62 => "01110", --   14
    63 => "01111", --   15
  );

  constant LUT_0_3_4_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11110", --   -2
    29 => "11110", --   -2
    30 => "11110", --   -2
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00011", --    3
    41 => "00100", --    4
    42 => "00101", --    5
    43 => "00110", --    6
    44 => "00111", --    7
    45 => "01000", --    8
    46 => "01001", --    9
    47 => "01001", --    9
    48 => "01010", --   10
    49 => "01010", --   10
    50 => "01010", --   10
    51 => "01011", --   11
    52 => "01011", --   11
    53 => "01011", --   11
    54 => "01100", --   12
    55 => "01100", --   12
    56 => "01100", --   12
    57 => "01101", --   13
    58 => "01101", --   13
    59 => "01101", --   13
    60 => "01110", --   14
    61 => "01110", --   14
    62 => "01110", --   14
    63 => "01111", --   15
  );

  constant LUT_0_3_5_DATA : lut_array_t_0 := (
    0 => "00100", --    4
    1 => "00101", --    5
    2 => "00101", --    5
    3 => "00110", --    6
    4 => "00111", --    7
    5 => "01000", --    8
    6 => "01001", --    9
    7 => "01001", --    9
    8 => "01010", --   10
    9 => "01010", --   10
    10 => "01011", --   11
    11 => "01011", --   11
    12 => "01011", --   11
    13 => "01011", --   11
    14 => "01011", --   11
    15 => "01011", --   11
    16 => "01011", --   11
    17 => "01010", --   10
    18 => "01010", --   10
    19 => "01010", --   10
    20 => "01001", --    9
    21 => "01001", --    9
    22 => "01000", --    8
    23 => "00111", --    7
    24 => "00111", --    7
    25 => "00110", --    6
    26 => "00100", --    4
    27 => "00011", --    3
    28 => "00010", --    2
    29 => "00000", --    0
    30 => "11110", --   -2
    31 => "11101", --   -3
    32 => "11100", --   -4
    33 => "11010", --   -6
    34 => "11001", --   -7
    35 => "11000", --   -8
    36 => "10111", --   -9
    37 => "10111", --   -9
    38 => "10110", --  -10
    39 => "10101", --  -11
    40 => "10100", --  -12
    41 => "10011", --  -13
    42 => "10010", --  -14
    43 => "10010", --  -14
    44 => "10001", --  -15
    45 => "10000", --  -16
    46 => "10000", --  -16
    47 => "10000", --  -16
    48 => "10000", --  -16
    49 => "10000", --  -16
    50 => "10000", --  -16
    51 => "10000", --  -16
    52 => "10000", --  -16
    53 => "10000", --  -16
    54 => "10000", --  -16
    55 => "10000", --  -16
    56 => "10000", --  -16
    57 => "10000", --  -16
    58 => "10000", --  -16
    59 => "10000", --  -16
    60 => "10000", --  -16
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_3_6_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11101", --   -3
    2 => "11101", --   -3
    3 => "11100", --   -4
    4 => "11011", --   -5
    5 => "11010", --   -6
    6 => "11001", --   -7
    7 => "11000", --   -8
    8 => "10111", --   -9
    9 => "10101", --  -11
    10 => "10100", --  -12
    11 => "10011", --  -13
    12 => "10010", --  -14
    13 => "10001", --  -15
    14 => "10000", --  -16
    15 => "10000", --  -16
    16 => "10000", --  -16
    17 => "10000", --  -16
    18 => "10000", --  -16
    19 => "10000", --  -16
    20 => "10000", --  -16
    21 => "10001", --  -15
    22 => "10010", --  -14
    23 => "10011", --  -13
    24 => "10100", --  -12
    25 => "10110", --  -10
    26 => "11000", --   -8
    27 => "11010", --   -6
    28 => "11100", --   -4
    29 => "11101", --   -3
    30 => "11111", --   -1
    31 => "00001", --    1
    32 => "00011", --    3
    33 => "00100", --    4
    34 => "00101", --    5
    35 => "00111", --    7
    36 => "01000", --    8
    37 => "01001", --    9
    38 => "01001", --    9
    39 => "01010", --   10
    40 => "01011", --   11
    41 => "01100", --   12
    42 => "01100", --   12
    43 => "01101", --   13
    44 => "01110", --   14
    45 => "01110", --   14
    46 => "01111", --   15
    47 => "01111", --   15
    48 => "01111", --   15
    49 => "01111", --   15
    50 => "01111", --   15
    51 => "01111", --   15
    52 => "01111", --   15
    53 => "01111", --   15
    54 => "01111", --   15
    55 => "01111", --   15
    56 => "01111", --   15
    57 => "01111", --   15
    58 => "01111", --   15
    59 => "01111", --   15
    60 => "01111", --   15
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_3_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11101", --   -3
    10 => "11101", --   -3
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11100", --   -4
    15 => "11100", --   -4
    16 => "11100", --   -4
    17 => "11101", --   -3
    18 => "11101", --   -3
    19 => "11101", --   -3
    20 => "11110", --   -2
    21 => "11111", --   -1
    22 => "00000", --    0
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00010", --    2
    26 => "00011", --    3
    27 => "00011", --    3
    28 => "00011", --    3
    29 => "00011", --    3
    30 => "00011", --    3
    31 => "00011", --    3
    32 => "00011", --    3
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00000", --    0
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11101", --   -3
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11100", --   -4
    50 => "11100", --   -4
    51 => "11100", --   -4
    52 => "11100", --   -4
    53 => "11100", --   -4
    54 => "11011", --   -5
    55 => "11011", --   -5
    56 => "11011", --   -5
    57 => "11010", --   -6
    58 => "11010", --   -6
    59 => "11001", --   -7
    60 => "11001", --   -7
    61 => "11000", --   -8
    62 => "11000", --   -8
    63 => "10111", --   -9
  );

  constant LUT_0_4_0_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00011", --    3
    8 => "00011", --    3
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00101", --    5
    12 => "00101", --    5
    13 => "00110", --    6
    14 => "00110", --    6
    15 => "00110", --    6
    16 => "00110", --    6
    17 => "00101", --    5
    18 => "00101", --    5
    19 => "00100", --    4
    20 => "00011", --    3
    21 => "00011", --    3
    22 => "00010", --    2
    23 => "00001", --    1
    24 => "00000", --    0
    25 => "11111", --   -1
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11110", --   -2
    29 => "11101", --   -3
    30 => "11101", --   -3
    31 => "11101", --   -3
    32 => "11101", --   -3
    33 => "11101", --   -3
    34 => "11101", --   -3
    35 => "11101", --   -3
    36 => "11101", --   -3
    37 => "11101", --   -3
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11100", --   -4
    43 => "11100", --   -4
    44 => "11100", --   -4
    45 => "11100", --   -4
    46 => "11100", --   -4
    47 => "11100", --   -4
    48 => "11100", --   -4
    49 => "11100", --   -4
    50 => "11011", --   -5
    51 => "11011", --   -5
    52 => "11011", --   -5
    53 => "11011", --   -5
    54 => "11010", --   -6
    55 => "11010", --   -6
    56 => "11010", --   -6
    57 => "11010", --   -6
    58 => "11001", --   -7
    59 => "11001", --   -7
    60 => "11001", --   -7
    61 => "11001", --   -7
    62 => "11001", --   -7
    63 => "11001", --   -7
  );

  constant LUT_0_4_1_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00011", --    3
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00101", --    5
    47 => "00101", --    5
    48 => "00101", --    5
    49 => "00110", --    6
    50 => "00110", --    6
    51 => "00110", --    6
    52 => "00110", --    6
    53 => "00110", --    6
    54 => "00110", --    6
    55 => "00110", --    6
    56 => "00110", --    6
    57 => "00110", --    6
    58 => "00110", --    6
    59 => "00110", --    6
    60 => "00110", --    6
    61 => "00110", --    6
    62 => "00110", --    6
    63 => "00110", --    6
  );

  constant LUT_0_4_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00011", --    3
    20 => "00011", --    3
    21 => "00011", --    3
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00010", --    2
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11100", --   -4
    41 => "11100", --   -4
    42 => "11100", --   -4
    43 => "11011", --   -5
    44 => "11011", --   -5
    45 => "11011", --   -5
    46 => "11011", --   -5
    47 => "11010", --   -6
    48 => "11010", --   -6
    49 => "11010", --   -6
    50 => "11010", --   -6
    51 => "11001", --   -7
    52 => "11001", --   -7
    53 => "11001", --   -7
    54 => "11000", --   -8
    55 => "11000", --   -8
    56 => "11000", --   -8
    57 => "10111", --   -9
    58 => "10111", --   -9
    59 => "10110", --  -10
    60 => "10110", --  -10
    61 => "10101", --  -11
    62 => "10101", --  -11
    63 => "10100", --  -12
  );

  constant LUT_0_4_3_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00011", --    3
    10 => "00011", --    3
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00011", --    3
    20 => "00011", --    3
    21 => "00011", --    3
    22 => "00011", --    3
    23 => "00010", --    2
    24 => "00010", --    2
    25 => "00010", --    2
    26 => "00010", --    2
    27 => "00010", --    2
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "11111", --   -1
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11100", --   -4
    41 => "11011", --   -5
    42 => "11011", --   -5
    43 => "11010", --   -6
    44 => "11001", --   -7
    45 => "11001", --   -7
    46 => "11000", --   -8
    47 => "10111", --   -9
    48 => "10111", --   -9
    49 => "10110", --  -10
    50 => "10110", --  -10
    51 => "10110", --  -10
    52 => "10110", --  -10
    53 => "10101", --  -11
    54 => "10101", --  -11
    55 => "10101", --  -11
    56 => "10101", --  -11
    57 => "10101", --  -11
    58 => "10101", --  -11
    59 => "10101", --  -11
    60 => "10101", --  -11
    61 => "10100", --  -12
    62 => "10100", --  -12
    63 => "10100", --  -12
  );

  constant LUT_0_4_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_4_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00011", --    3
    42 => "00011", --    3
    43 => "00100", --    4
    44 => "00100", --    4
    45 => "00101", --    5
    46 => "00101", --    5
    47 => "00110", --    6
    48 => "00110", --    6
    49 => "00110", --    6
    50 => "00111", --    7
    51 => "00111", --    7
    52 => "00111", --    7
    53 => "00111", --    7
    54 => "01000", --    8
    55 => "01000", --    8
    56 => "01000", --    8
    57 => "01001", --    9
    58 => "01001", --    9
    59 => "01001", --    9
    60 => "01010", --   10
    61 => "01010", --   10
    62 => "01011", --   11
    63 => "01011", --   11
  );

  constant LUT_0_4_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11101", --   -3
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11100", --   -4
    14 => "11100", --   -4
    15 => "11100", --   -4
    16 => "11100", --   -4
    17 => "11101", --   -3
    18 => "11101", --   -3
    19 => "11101", --   -3
    20 => "11101", --   -3
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00010", --    2
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00100", --    4
    60 => "00101", --    5
    61 => "00101", --    5
    62 => "00101", --    5
    63 => "00110", --    6
  );

  constant LUT_0_4_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11110", --   -2
    14 => "11110", --   -2
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00011", --    3
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00100", --    4
    51 => "00100", --    4
    52 => "00101", --    5
    53 => "00101", --    5
    54 => "00101", --    5
    55 => "00110", --    6
    56 => "00110", --    6
    57 => "00111", --    7
    58 => "00111", --    7
    59 => "01000", --    8
    60 => "01000", --    8
    61 => "01000", --    8
    62 => "01000", --    8
    63 => "01000", --    8
  );

  constant LUT_0_5_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "00000", --    0
    54 => "00000", --    0
    55 => "00000", --    0
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "00000", --    0
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_5_1_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00100", --    4
    45 => "00100", --    4
    46 => "00100", --    4
    47 => "00101", --    5
    48 => "00101", --    5
    49 => "00101", --    5
    50 => "00101", --    5
    51 => "00101", --    5
    52 => "00110", --    6
    53 => "00110", --    6
    54 => "00110", --    6
    55 => "00110", --    6
    56 => "00110", --    6
    57 => "00110", --    6
    58 => "00111", --    7
    59 => "00111", --    7
    60 => "00111", --    7
    61 => "00111", --    7
    62 => "00111", --    7
    63 => "01000", --    8
  );

  constant LUT_0_5_2_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_5_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00001", --    1
    57 => "00001", --    1
    58 => "00001", --    1
    59 => "00001", --    1
    60 => "00001", --    1
    61 => "00001", --    1
    62 => "00001", --    1
    63 => "00001", --    1
  );

  constant LUT_0_5_4_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11101", --   -3
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11101", --   -3
    19 => "11101", --   -3
    20 => "11101", --   -3
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00010", --    2
    32 => "00010", --    2
    33 => "00010", --    2
    34 => "00011", --    3
    35 => "00011", --    3
    36 => "00011", --    3
    37 => "00100", --    4
    38 => "00100", --    4
    39 => "00101", --    5
    40 => "00101", --    5
    41 => "00110", --    6
    42 => "00110", --    6
    43 => "00111", --    7
    44 => "00111", --    7
    45 => "01000", --    8
    46 => "01000", --    8
    47 => "01001", --    9
    48 => "01010", --   10
    49 => "01010", --   10
    50 => "01011", --   11
    51 => "01011", --   11
    52 => "01100", --   12
    53 => "01100", --   12
    54 => "01101", --   13
    55 => "01101", --   13
    56 => "01110", --   14
    57 => "01111", --   15
    58 => "01111", --   15
    59 => "01111", --   15
    60 => "01111", --   15
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_5_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11101", --   -3
    5 => "11100", --   -4
    6 => "11010", --   -6
    7 => "11001", --   -7
    8 => "10111", --   -9
    9 => "10110", --  -10
    10 => "10101", --  -11
    11 => "10100", --  -12
    12 => "10011", --  -13
    13 => "10100", --  -12
    14 => "10100", --  -12
    15 => "10110", --  -10
    16 => "10111", --   -9
    17 => "11001", --   -7
    18 => "11011", --   -5
    19 => "11101", --   -3
    20 => "11110", --   -2
    21 => "00000", --    0
    22 => "00001", --    1
    23 => "00010", --    2
    24 => "00011", --    3
    25 => "00011", --    3
    26 => "00100", --    4
    27 => "00100", --    4
    28 => "00100", --    4
    29 => "00011", --    3
    30 => "00011", --    3
    31 => "00011", --    3
    32 => "00010", --    2
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00010", --    2
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_5_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00011", --    3
    45 => "00011", --    3
    46 => "00011", --    3
    47 => "00100", --    4
    48 => "00100", --    4
    49 => "00100", --    4
    50 => "00100", --    4
    51 => "00100", --    4
    52 => "00101", --    5
    53 => "00101", --    5
    54 => "00101", --    5
    55 => "00101", --    5
    56 => "00101", --    5
    57 => "00110", --    6
    58 => "00110", --    6
    59 => "00110", --    6
    60 => "00110", --    6
    61 => "00111", --    7
    62 => "00111", --    7
    63 => "00111", --    7
  );

  constant LUT_0_5_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00011", --    3
    45 => "00100", --    4
    46 => "00100", --    4
    47 => "00100", --    4
    48 => "00101", --    5
    49 => "00101", --    5
    50 => "00101", --    5
    51 => "00110", --    6
    52 => "00110", --    6
    53 => "00111", --    7
    54 => "00111", --    7
    55 => "00111", --    7
    56 => "01000", --    8
    57 => "01000", --    8
    58 => "01000", --    8
    59 => "01001", --    9
    60 => "01001", --    9
    61 => "01001", --    9
    62 => "01001", --    9
    63 => "01001", --    9
  );

  constant LUT_0_6_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "00000", --    0
    54 => "00000", --    0
    55 => "00000", --    0
    56 => "00000", --    0
    57 => "00000", --    0
    58 => "00000", --    0
    59 => "00000", --    0
    60 => "00000", --    0
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_6_1_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_6_2_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_6_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_6_4_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11110", --   -2
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11100", --   -4
    53 => "11100", --   -4
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11100", --   -4
    57 => "11011", --   -5
    58 => "11011", --   -5
    59 => "11011", --   -5
    60 => "11010", --   -6
    61 => "11010", --   -6
    62 => "11010", --   -6
    63 => "11001", --   -7
  );

  constant LUT_0_6_5_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_6_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "00000", --    0
    54 => "00000", --    0
    55 => "00001", --    1
    56 => "00001", --    1
    57 => "00001", --    1
    58 => "00001", --    1
    59 => "00001", --    1
    60 => "00001", --    1
    61 => "00001", --    1
    62 => "00001", --    1
    63 => "00001", --    1
  );

  constant LUT_0_6_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_7_0_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11101", --   -3
    7 => "11101", --   -3
    8 => "11101", --   -3
    9 => "11101", --   -3
    10 => "11100", --   -4
    11 => "11100", --   -4
    12 => "11100", --   -4
    13 => "11100", --   -4
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00011", --    3
    47 => "00011", --    3
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00100", --    4
    54 => "00100", --    4
    55 => "00100", --    4
    56 => "00100", --    4
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00100", --    4
    60 => "00101", --    5
    61 => "00101", --    5
    62 => "00101", --    5
    63 => "00101", --    5
  );

  constant LUT_0_7_1_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_7_2_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11110", --   -2
    14 => "11110", --   -2
    15 => "11110", --   -2
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_7_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11110", --   -2
    14 => "11110", --   -2
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11110", --   -2
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00011", --    3
    45 => "00011", --    3
    46 => "00011", --    3
    47 => "00011", --    3
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00100", --    4
    55 => "00100", --    4
    56 => "00100", --    4
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00100", --    4
    60 => "00100", --    4
    61 => "00100", --    4
    62 => "00101", --    5
    63 => "00101", --    5
  );

  constant LUT_0_7_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11110", --   -2
    14 => "11110", --   -2
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11110", --   -2
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00100", --    4
    62 => "00100", --    4
    63 => "00100", --    4
  );

  constant LUT_0_7_5_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00010", --    2
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00011", --    3
    5 => "00011", --    3
    6 => "00011", --    3
    7 => "00011", --    3
    8 => "00100", --    4
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11110", --   -2
    29 => "11110", --   -2
    30 => "11110", --   -2
    31 => "11101", --   -3
    32 => "11101", --   -3
    33 => "11101", --   -3
    34 => "11110", --   -2
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11110", --   -2
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_7_6_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11101", --   -3
    10 => "11101", --   -3
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11110", --   -2
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11110", --   -2
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00010", --    2
    29 => "00010", --    2
    30 => "00010", --    2
    31 => "00010", --    2
    32 => "00010", --    2
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00010", --    2
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00011", --    3
    49 => "00011", --    3
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_7_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00010", --    2
    63 => "00011", --    3
  );

  constant LUT_0_8_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11110", --   -2
  );

  constant LUT_0_8_1_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_8_2_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_8_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11110", --   -2
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11100", --   -4
    57 => "11100", --   -4
    58 => "11100", --   -4
    59 => "11011", --   -5
    60 => "11011", --   -5
    61 => "11011", --   -5
    62 => "11011", --   -5
    63 => "11011", --   -5
  );

  constant LUT_0_8_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_8_5_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00010", --    2
    63 => "00010", --    2
  );

  constant LUT_0_8_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11101", --   -3
  );

  constant LUT_0_8_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11111", --   -1
  );

  constant LUT_0_9_0_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00100", --    4
    63 => "00100", --    4
  );

  constant LUT_0_9_1_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_9_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_9_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11110", --   -2
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11100", --   -4
    53 => "11100", --   -4
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11100", --   -4
    57 => "11011", --   -5
    58 => "11011", --   -5
    59 => "11011", --   -5
    60 => "11011", --   -5
    61 => "11010", --   -6
    62 => "11010", --   -6
    63 => "11010", --   -6
  );

  constant LUT_0_9_4_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00010", --    2
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00011", --    3
    44 => "00011", --    3
    45 => "00011", --    3
    46 => "00100", --    4
    47 => "00100", --    4
    48 => "00100", --    4
    49 => "00101", --    5
    50 => "00101", --    5
    51 => "00101", --    5
    52 => "00110", --    6
    53 => "00110", --    6
    54 => "00110", --    6
    55 => "00111", --    7
    56 => "00111", --    7
    57 => "00111", --    7
    58 => "01000", --    8
    59 => "01000", --    8
    60 => "01001", --    9
    61 => "01001", --    9
    62 => "01001", --    9
    63 => "01010", --   10
  );

  constant LUT_0_9_5_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11100", --   -4
    57 => "11100", --   -4
    58 => "11100", --   -4
    59 => "11100", --   -4
    60 => "11100", --   -4
    61 => "11011", --   -5
    62 => "11011", --   -5
    63 => "11011", --   -5
  );

  constant LUT_0_9_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_9_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00010", --    2
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00100", --    4
    60 => "00100", --    4
    61 => "00100", --    4
    62 => "00101", --    5
    63 => "00101", --    5
  );

  constant LUT_0_10_0_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_10_1_DATA : lut_array_t_0 := (
    0 => "11011", --   -5
    1 => "11011", --   -5
    2 => "11011", --   -5
    3 => "11010", --   -6
    4 => "11010", --   -6
    5 => "11010", --   -6
    6 => "11010", --   -6
    7 => "11010", --   -6
    8 => "11010", --   -6
    9 => "11010", --   -6
    10 => "11011", --   -5
    11 => "11011", --   -5
    12 => "11011", --   -5
    13 => "11100", --   -4
    14 => "11100", --   -4
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00010", --    2
    36 => "00011", --    3
    37 => "00011", --    3
    38 => "00011", --    3
    39 => "00100", --    4
    40 => "00100", --    4
    41 => "00100", --    4
    42 => "00100", --    4
    43 => "00101", --    5
    44 => "00101", --    5
    45 => "00101", --    5
    46 => "00101", --    5
    47 => "00110", --    6
    48 => "00110", --    6
    49 => "00110", --    6
    50 => "00111", --    7
    51 => "00111", --    7
    52 => "00111", --    7
    53 => "01000", --    8
    54 => "01000", --    8
    55 => "01001", --    9
    56 => "01001", --    9
    57 => "01001", --    9
    58 => "01010", --   10
    59 => "01010", --   10
    60 => "01011", --   11
    61 => "01011", --   11
    62 => "01011", --   11
    63 => "01100", --   12
  );

  constant LUT_0_10_2_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00010", --    2
    63 => "00010", --    2
  );

  constant LUT_0_10_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11110", --   -2
    41 => "11101", --   -3
    42 => "11101", --   -3
    43 => "11101", --   -3
    44 => "11100", --   -4
    45 => "11100", --   -4
    46 => "11100", --   -4
    47 => "11100", --   -4
    48 => "11011", --   -5
    49 => "11011", --   -5
    50 => "11011", --   -5
    51 => "11011", --   -5
    52 => "11010", --   -6
    53 => "11010", --   -6
    54 => "11010", --   -6
    55 => "11001", --   -7
    56 => "11001", --   -7
    57 => "11001", --   -7
    58 => "11000", --   -8
    59 => "11000", --   -8
    60 => "11000", --   -8
    61 => "10111", --   -9
    62 => "10111", --   -9
    63 => "10110", --  -10
  );

  constant LUT_0_10_4_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00010", --    2
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00011", --    3
    51 => "00011", --    3
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00100", --    4
    56 => "00100", --    4
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00101", --    5
    60 => "00101", --    5
    61 => "00101", --    5
    62 => "00101", --    5
    63 => "00101", --    5
  );

  constant LUT_0_10_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00001", --    1
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00100", --    4
    62 => "00100", --    4
    63 => "00100", --    4
  );

  constant LUT_0_10_6_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00010", --    2
    2 => "00010", --    2
    3 => "00011", --    3
    4 => "00011", --    3
    5 => "00100", --    4
    6 => "00100", --    4
    7 => "00100", --    4
    8 => "00100", --    4
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00100", --    4
    12 => "00100", --    4
    13 => "00100", --    4
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11110", --   -2
    34 => "11110", --   -2
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11101", --   -3
    57 => "11100", --   -4
    58 => "11100", --   -4
    59 => "11100", --   -4
    60 => "11011", --   -5
    61 => "11011", --   -5
    62 => "11011", --   -5
    63 => "11010", --   -6
  );

  constant LUT_0_10_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11101", --   -3
  );

  constant LUT_0_11_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "00000", --    0
    54 => "00000", --    0
    55 => "00000", --    0
    56 => "00000", --    0
    57 => "00000", --    0
    58 => "00000", --    0
    59 => "00000", --    0
    60 => "00001", --    1
    61 => "00001", --    1
    62 => "00001", --    1
    63 => "00000", --    0
  );

  constant LUT_0_11_1_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11101", --   -3
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11100", --   -4
    43 => "11100", --   -4
    44 => "11100", --   -4
    45 => "11100", --   -4
    46 => "11011", --   -5
    47 => "11011", --   -5
    48 => "11011", --   -5
    49 => "11010", --   -6
    50 => "11010", --   -6
    51 => "11001", --   -7
    52 => "11001", --   -7
    53 => "11001", --   -7
    54 => "11000", --   -8
    55 => "11000", --   -8
    56 => "10111", --   -9
    57 => "10111", --   -9
    58 => "10111", --   -9
    59 => "10110", --  -10
    60 => "10110", --  -10
    61 => "10101", --  -11
    62 => "10101", --  -11
    63 => "10101", --  -11
  );

  constant LUT_0_11_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00011", --    3
    9 => "00011", --    3
    10 => "00011", --    3
    11 => "00011", --    3
    12 => "00011", --    3
    13 => "00011", --    3
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11100", --   -4
    57 => "11100", --   -4
    58 => "11100", --   -4
    59 => "11100", --   -4
    60 => "11100", --   -4
    61 => "11100", --   -4
    62 => "11100", --   -4
    63 => "11100", --   -4
  );

  constant LUT_0_11_3_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00011", --    3
    5 => "00011", --    3
    6 => "00011", --    3
    7 => "00100", --    4
    8 => "00100", --    4
    9 => "00100", --    4
    10 => "00101", --    5
    11 => "00101", --    5
    12 => "00101", --    5
    13 => "00101", --    5
    14 => "00101", --    5
    15 => "00101", --    5
    16 => "00100", --    4
    17 => "00100", --    4
    18 => "00100", --    4
    19 => "00011", --    3
    20 => "00011", --    3
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11110", --   -2
    33 => "11110", --   -2
    34 => "11110", --   -2
    35 => "11110", --   -2
    36 => "11101", --   -3
    37 => "11101", --   -3
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11101", --   -3
    43 => "11101", --   -3
    44 => "11101", --   -3
    45 => "11100", --   -4
    46 => "11100", --   -4
    47 => "11100", --   -4
    48 => "11100", --   -4
    49 => "11100", --   -4
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11101", --   -3
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_11_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00100", --    4
    58 => "00100", --    4
    59 => "00100", --    4
    60 => "00100", --    4
    61 => "00101", --    5
    62 => "00101", --    5
    63 => "00101", --    5
  );

  constant LUT_0_11_5_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11101", --   -3
    57 => "11101", --   -3
    58 => "11101", --   -3
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11100", --   -4
    63 => "11100", --   -4
  );

  constant LUT_0_11_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11101", --   -3
  );

  constant LUT_0_11_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11101", --   -3
    9 => "11101", --   -3
    10 => "11101", --   -3
    11 => "11101", --   -3
    12 => "11101", --   -3
    13 => "11101", --   -3
    14 => "11101", --   -3
    15 => "11101", --   -3
    16 => "11101", --   -3
    17 => "11101", --   -3
    18 => "11101", --   -3
    19 => "11101", --   -3
    20 => "11101", --   -3
    21 => "11101", --   -3
    22 => "11101", --   -3
    23 => "11101", --   -3
    24 => "11101", --   -3
    25 => "11101", --   -3
    26 => "11110", --   -2
    27 => "11110", --   -2
    28 => "11110", --   -2
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00001", --    1
    34 => "00001", --    1
    35 => "00010", --    2
    36 => "00010", --    2
    37 => "00010", --    2
    38 => "00011", --    3
    39 => "00011", --    3
    40 => "00100", --    4
    41 => "00100", --    4
    42 => "00101", --    5
    43 => "00101", --    5
    44 => "00110", --    6
    45 => "00110", --    6
    46 => "00110", --    6
    47 => "00111", --    7
    48 => "00111", --    7
    49 => "01000", --    8
    50 => "01000", --    8
    51 => "01000", --    8
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01010", --   10
    57 => "01011", --   11
    58 => "01011", --   11
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01101", --   13
    62 => "01101", --   13
    63 => "01101", --   13
  );

  constant LUT_0_12_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11101", --   -3
    56 => "11101", --   -3
    57 => "11101", --   -3
    58 => "11101", --   -3
    59 => "11100", --   -4
    60 => "11100", --   -4
    61 => "11100", --   -4
    62 => "11100", --   -4
    63 => "11100", --   -4
  );

  constant LUT_0_12_1_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00010", --    2
    46 => "00010", --    2
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00011", --    3
    53 => "00011", --    3
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_12_2_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11111", --   -1
    48 => "11111", --   -1
    49 => "11111", --   -1
    50 => "11111", --   -1
    51 => "11111", --   -1
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_12_3_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_12_4_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00010", --    2
    55 => "00010", --    2
    56 => "00010", --    2
    57 => "00010", --    2
    58 => "00010", --    2
    59 => "00011", --    3
    60 => "00011", --    3
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_12_5_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "11111", --   -1
    17 => "11111", --   -1
    18 => "11111", --   -1
    19 => "11111", --   -1
    20 => "11111", --   -1
    21 => "11111", --   -1
    22 => "11111", --   -1
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00001", --    1
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00010", --    2
    43 => "00011", --    3
    44 => "00011", --    3
    45 => "00011", --    3
    46 => "00011", --    3
    47 => "00100", --    4
    48 => "00100", --    4
    49 => "00100", --    4
    50 => "00101", --    5
    51 => "00101", --    5
    52 => "00101", --    5
    53 => "00101", --    5
    54 => "00110", --    6
    55 => "00110", --    6
    56 => "00110", --    6
    57 => "00111", --    7
    58 => "00111", --    7
    59 => "00111", --    7
    60 => "01000", --    8
    61 => "01000", --    8
    62 => "01000", --    8
    63 => "01001", --    9
  );

  constant LUT_0_12_6_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11110", --   -2
    41 => "11110", --   -2
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11101", --   -3
    45 => "11101", --   -3
    46 => "11101", --   -3
    47 => "11101", --   -3
    48 => "11101", --   -3
    49 => "11101", --   -3
    50 => "11100", --   -4
    51 => "11100", --   -4
    52 => "11100", --   -4
    53 => "11100", --   -4
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11011", --   -5
    57 => "11011", --   -5
    58 => "11011", --   -5
    59 => "11011", --   -5
    60 => "11010", --   -6
    61 => "11010", --   -6
    62 => "11010", --   -6
    63 => "11010", --   -6
  );

  constant LUT_0_12_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00010", --    2
    17 => "00010", --    2
    18 => "00010", --    2
    19 => "00010", --    2
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00010", --    2
    25 => "00010", --    2
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11110", --   -2
    38 => "11110", --   -2
    39 => "11110", --   -2
    40 => "11101", --   -3
    41 => "11101", --   -3
    42 => "11100", --   -4
    43 => "11100", --   -4
    44 => "11011", --   -5
    45 => "11011", --   -5
    46 => "11010", --   -6
    47 => "11010", --   -6
    48 => "11001", --   -7
    49 => "11001", --   -7
    50 => "11000", --   -8
    51 => "11000", --   -8
    52 => "10111", --   -9
    53 => "10111", --   -9
    54 => "10110", --  -10
    55 => "10110", --  -10
    56 => "10101", --  -11
    57 => "10101", --  -11
    58 => "10100", --  -12
    59 => "10100", --  -12
    60 => "10011", --  -13
    61 => "10011", --  -13
    62 => "10010", --  -14
    63 => "10010", --  -14
  );

  constant LUT_0_13_0_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "00000", --    0
    53 => "00000", --    0
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11111", --   -1
    61 => "11111", --   -1
    62 => "11111", --   -1
    63 => "11110", --   -2
  );

  constant LUT_0_13_1_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11110", --   -2
    43 => "11110", --   -2
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11101", --   -3
    59 => "11101", --   -3
    60 => "11101", --   -3
    61 => "11101", --   -3
    62 => "11101", --   -3
    63 => "11101", --   -3
  );

  constant LUT_0_13_2_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00000", --    0
    43 => "00000", --    0
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00001", --    1
    57 => "00001", --    1
    58 => "00001", --    1
    59 => "00001", --    1
    60 => "00001", --    1
    61 => "00000", --    0
    62 => "00000", --    0
    63 => "00000", --    0
  );

  constant LUT_0_13_3_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "00000", --    0
    11 => "00000", --    0
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00001", --    1
    40 => "00001", --    1
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00010", --    2
    48 => "00010", --    2
    49 => "00010", --    2
    50 => "00010", --    2
    51 => "00010", --    2
    52 => "00010", --    2
    53 => "00010", --    2
    54 => "00011", --    3
    55 => "00011", --    3
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00011", --    3
    59 => "00011", --    3
    60 => "00100", --    4
    61 => "00100", --    4
    62 => "00100", --    4
    63 => "00100", --    4
  );

  constant LUT_0_13_4_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00001", --    1
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11110", --   -2
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11101", --   -3
    55 => "11101", --   -3
    56 => "11100", --   -4
    57 => "11100", --   -4
    58 => "11100", --   -4
    59 => "11100", --   -4
    60 => "11011", --   -5
    61 => "11011", --   -5
    62 => "11011", --   -5
    63 => "11011", --   -5
  );

  constant LUT_0_13_5_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00001", --    1
    2 => "00001", --    1
    3 => "00010", --    2
    4 => "00010", --    2
    5 => "00010", --    2
    6 => "00010", --    2
    7 => "00010", --    2
    8 => "00010", --    2
    9 => "00010", --    2
    10 => "00010", --    2
    11 => "00010", --    2
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00010", --    2
    15 => "00010", --    2
    16 => "00010", --    2
    17 => "00001", --    1
    18 => "00001", --    1
    19 => "00001", --    1
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "11111", --   -1
    39 => "11111", --   -1
    40 => "11111", --   -1
    41 => "11111", --   -1
    42 => "11111", --   -1
    43 => "11111", --   -1
    44 => "11111", --   -1
    45 => "11110", --   -2
    46 => "11110", --   -2
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "11110", --   -2
    53 => "11110", --   -2
    54 => "11110", --   -2
    55 => "11110", --   -2
    56 => "11110", --   -2
    57 => "11110", --   -2
    58 => "11110", --   -2
    59 => "11110", --   -2
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_13_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00000", --    0
    5 => "00000", --    0
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00000", --    0
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "00000", --    0
    13 => "00000", --    0
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "00000", --    0
    24 => "00000", --    0
    25 => "00000", --    0
    26 => "00000", --    0
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00001", --    1
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00001", --    1
    45 => "00001", --    1
    46 => "00001", --    1
    47 => "00001", --    1
    48 => "00001", --    1
    49 => "00001", --    1
    50 => "00001", --    1
    51 => "00001", --    1
    52 => "00001", --    1
    53 => "00001", --    1
    54 => "00001", --    1
    55 => "00001", --    1
    56 => "00001", --    1
    57 => "00001", --    1
    58 => "00001", --    1
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00010", --    2
    62 => "00010", --    2
    63 => "00010", --    2
  );

  constant LUT_0_13_7_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "00000", --    0
    2 => "00000", --    0
    3 => "00000", --    0
    4 => "00001", --    1
    5 => "00001", --    1
    6 => "00001", --    1
    7 => "00001", --    1
    8 => "00001", --    1
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00001", --    1
    13 => "00001", --    1
    14 => "00001", --    1
    15 => "00001", --    1
    16 => "00001", --    1
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11111", --   -1
    32 => "11111", --   -1
    33 => "00000", --    0
    34 => "00000", --    0
    35 => "00000", --    0
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00000", --    0
    39 => "00000", --    0
    40 => "00000", --    0
    41 => "00000", --    0
    42 => "00001", --    1
    43 => "00001", --    1
    44 => "00000", --    0
    45 => "00000", --    0
    46 => "00000", --    0
    47 => "00000", --    0
    48 => "00000", --    0
    49 => "00000", --    0
    50 => "00000", --    0
    51 => "00000", --    0
    52 => "11111", --   -1
    53 => "11111", --   -1
    54 => "11111", --   -1
    55 => "11111", --   -1
    56 => "11111", --   -1
    57 => "11111", --   -1
    58 => "11111", --   -1
    59 => "11111", --   -1
    60 => "11110", --   -2
    61 => "11110", --   -2
    62 => "11110", --   -2
    63 => "11110", --   -2
  );

  constant LUT_0_14_0_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11110", --   -2
    9 => "11110", --   -2
    10 => "11110", --   -2
    11 => "11110", --   -2
    12 => "11110", --   -2
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00001", --    1
    21 => "00001", --    1
    22 => "00001", --    1
    23 => "00001", --    1
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "11110", --   -2
    32 => "11110", --   -2
    33 => "11110", --   -2
    34 => "11110", --   -2
    35 => "11110", --   -2
    36 => "11111", --   -1
    37 => "11111", --   -1
    38 => "00000", --    0
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00010", --    2
    42 => "00011", --    3
    43 => "00100", --    4
    44 => "00101", --    5
    45 => "00101", --    5
    46 => "00110", --    6
    47 => "00111", --    7
    48 => "00111", --    7
    49 => "01000", --    8
    50 => "01000", --    8
    51 => "01001", --    9
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01011", --   11
    57 => "01011", --   11
    58 => "01100", --   12
    59 => "01100", --   12
    60 => "01101", --   13
    61 => "01110", --   14
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_14_1_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11110", --   -2
    7 => "11110", --   -2
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "00000", --    0
    15 => "00000", --    0
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00000", --    0
    19 => "00000", --    0
    20 => "00000", --    0
    21 => "00000", --    0
    22 => "00000", --    0
    23 => "11111", --   -1
    24 => "11111", --   -1
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11110", --   -2
    30 => "11110", --   -2
    31 => "11110", --   -2
    32 => "11110", --   -2
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11111", --   -1
    36 => "00000", --    0
    37 => "00000", --    0
    38 => "00001", --    1
    39 => "00001", --    1
    40 => "00010", --    2
    41 => "00011", --    3
    42 => "00011", --    3
    43 => "00100", --    4
    44 => "00100", --    4
    45 => "00101", --    5
    46 => "00101", --    5
    47 => "00101", --    5
    48 => "00101", --    5
    49 => "00101", --    5
    50 => "00101", --    5
    51 => "00101", --    5
    52 => "00101", --    5
    53 => "00100", --    4
    54 => "00100", --    4
    55 => "00100", --    4
    56 => "00011", --    3
    57 => "00011", --    3
    58 => "00010", --    2
    59 => "00010", --    2
    60 => "00010", --    2
    61 => "00011", --    3
    62 => "00011", --    3
    63 => "00011", --    3
  );

  constant LUT_0_14_2_DATA : lut_array_t_0 := (
    0 => "11100", --   -4
    1 => "11100", --   -4
    2 => "11011", --   -5
    3 => "11011", --   -5
    4 => "11011", --   -5
    5 => "11011", --   -5
    6 => "11011", --   -5
    7 => "11011", --   -5
    8 => "11010", --   -6
    9 => "11010", --   -6
    10 => "11010", --   -6
    11 => "11010", --   -6
    12 => "11010", --   -6
    13 => "11001", --   -7
    14 => "11001", --   -7
    15 => "11000", --   -8
    16 => "10111", --   -9
    17 => "10111", --   -9
    18 => "10111", --   -9
    19 => "10111", --   -9
    20 => "10111", --   -9
    21 => "10111", --   -9
    22 => "10111", --   -9
    23 => "11000", --   -8
    24 => "11000", --   -8
    25 => "11001", --   -7
    26 => "11010", --   -6
    27 => "11011", --   -5
    28 => "11100", --   -4
    29 => "11101", --   -3
    30 => "11110", --   -2
    31 => "11111", --   -1
    32 => "00001", --    1
    33 => "00010", --    2
    34 => "00011", --    3
    35 => "00100", --    4
    36 => "00110", --    6
    37 => "00111", --    7
    38 => "00111", --    7
    39 => "01000", --    8
    40 => "01000", --    8
    41 => "01000", --    8
    42 => "01000", --    8
    43 => "01000", --    8
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "00111", --    7
    47 => "00111", --    7
    48 => "00111", --    7
    49 => "01000", --    8
    50 => "01000", --    8
    51 => "01000", --    8
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01001", --    9
    55 => "01001", --    9
    56 => "01010", --   10
    57 => "01010", --   10
    58 => "01011", --   11
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01101", --   13
    62 => "01110", --   14
    63 => "01111", --   15
  );

  constant LUT_0_14_3_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "00000", --    0
    7 => "00000", --    0
    8 => "00000", --    0
    9 => "00001", --    1
    10 => "00001", --    1
    11 => "00001", --    1
    12 => "00010", --    2
    13 => "00010", --    2
    14 => "00011", --    3
    15 => "00011", --    3
    16 => "00011", --    3
    17 => "00100", --    4
    18 => "00100", --    4
    19 => "00101", --    5
    20 => "00110", --    6
    21 => "00110", --    6
    22 => "00111", --    7
    23 => "00111", --    7
    24 => "01000", --    8
    25 => "01000", --    8
    26 => "01000", --    8
    27 => "01000", --    8
    28 => "00111", --    7
    29 => "00111", --    7
    30 => "00110", --    6
    31 => "00100", --    4
    32 => "00011", --    3
    33 => "00001", --    1
    34 => "11111", --   -1
    35 => "11110", --   -2
    36 => "11100", --   -4
    37 => "11011", --   -5
    38 => "11001", --   -7
    39 => "11001", --   -7
    40 => "11000", --   -8
    41 => "11000", --   -8
    42 => "11001", --   -7
    43 => "11001", --   -7
    44 => "11010", --   -6
    45 => "11011", --   -5
    46 => "11011", --   -5
    47 => "11100", --   -4
    48 => "11100", --   -4
    49 => "11101", --   -3
    50 => "11110", --   -2
    51 => "11110", --   -2
    52 => "00000", --    0
    53 => "00001", --    1
    54 => "00010", --    2
    55 => "00100", --    4
    56 => "00101", --    5
    57 => "00110", --    6
    58 => "00111", --    7
    59 => "00111", --    7
    60 => "00110", --    6
    61 => "00101", --    5
    62 => "00100", --    4
    63 => "00011", --    3
  );

  constant LUT_0_14_4_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11101", --   -3
    2 => "11101", --   -3
    3 => "11101", --   -3
    4 => "11101", --   -3
    5 => "11101", --   -3
    6 => "11101", --   -3
    7 => "11101", --   -3
    8 => "11101", --   -3
    9 => "11101", --   -3
    10 => "11101", --   -3
    11 => "11101", --   -3
    12 => "11110", --   -2
    13 => "11110", --   -2
    14 => "11111", --   -1
    15 => "11111", --   -1
    16 => "00000", --    0
    17 => "00000", --    0
    18 => "00001", --    1
    19 => "00010", --    2
    20 => "00011", --    3
    21 => "00100", --    4
    22 => "00101", --    5
    23 => "00110", --    6
    24 => "00111", --    7
    25 => "00111", --    7
    26 => "00111", --    7
    27 => "00111", --    7
    28 => "00110", --    6
    29 => "00101", --    5
    30 => "00100", --    4
    31 => "00011", --    3
    32 => "00001", --    1
    33 => "00000", --    0
    34 => "11110", --   -2
    35 => "11101", --   -3
    36 => "11100", --   -4
    37 => "11011", --   -5
    38 => "11011", --   -5
    39 => "11011", --   -5
    40 => "11100", --   -4
    41 => "11110", --   -2
    42 => "00000", --    0
    43 => "00010", --    2
    44 => "00100", --    4
    45 => "00111", --    7
    46 => "01001", --    9
    47 => "01100", --   12
    48 => "01110", --   14
    49 => "01111", --   15
    50 => "01111", --   15
    51 => "01111", --   15
    52 => "01111", --   15
    53 => "01111", --   15
    54 => "01111", --   15
    55 => "01111", --   15
    56 => "01111", --   15
    57 => "01111", --   15
    58 => "01110", --   14
    59 => "01101", --   13
    60 => "01100", --   12
    61 => "01011", --   11
    62 => "01011", --   11
    63 => "01010", --   10
  );

  constant LUT_0_14_5_DATA : lut_array_t_0 := (
    0 => "00111", --    7
    1 => "01000", --    8
    2 => "01001", --    9
    3 => "01010", --   10
    4 => "01011", --   11
    5 => "01011", --   11
    6 => "01100", --   12
    7 => "01100", --   12
    8 => "01100", --   12
    9 => "01100", --   12
    10 => "01100", --   12
    11 => "01100", --   12
    12 => "01011", --   11
    13 => "01011", --   11
    14 => "01010", --   10
    15 => "01010", --   10
    16 => "01001", --    9
    17 => "01000", --    8
    18 => "01000", --    8
    19 => "00111", --    7
    20 => "00111", --    7
    21 => "00111", --    7
    22 => "00111", --    7
    23 => "00111", --    7
    24 => "00111", --    7
    25 => "00110", --    6
    26 => "00110", --    6
    27 => "00101", --    5
    28 => "00100", --    4
    29 => "00011", --    3
    30 => "00010", --    2
    31 => "00001", --    1
    32 => "00000", --    0
    33 => "11111", --   -1
    34 => "11101", --   -3
    35 => "11100", --   -4
    36 => "11011", --   -5
    37 => "11010", --   -6
    38 => "11001", --   -7
    39 => "11000", --   -8
    40 => "11000", --   -8
    41 => "10111", --   -9
    42 => "10111", --   -9
    43 => "10110", --  -10
    44 => "10101", --  -11
    45 => "10100", --  -12
    46 => "10011", --  -13
    47 => "10010", --  -14
    48 => "10001", --  -15
    49 => "10000", --  -16
    50 => "10000", --  -16
    51 => "10000", --  -16
    52 => "10000", --  -16
    53 => "10000", --  -16
    54 => "10000", --  -16
    55 => "10000", --  -16
    56 => "10000", --  -16
    57 => "10000", --  -16
    58 => "10000", --  -16
    59 => "10000", --  -16
    60 => "10000", --  -16
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_14_6_DATA : lut_array_t_0 := (
    0 => "00000", --    0
    1 => "11111", --   -1
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11101", --   -3
    5 => "11101", --   -3
    6 => "11100", --   -4
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11101", --   -3
    12 => "11110", --   -2
    13 => "11111", --   -1
    14 => "00001", --    1
    15 => "00011", --    3
    16 => "00101", --    5
    17 => "01000", --    8
    18 => "01010", --   10
    19 => "01100", --   12
    20 => "01110", --   14
    21 => "01111", --   15
    22 => "01111", --   15
    23 => "01111", --   15
    24 => "01111", --   15
    25 => "01111", --   15
    26 => "01111", --   15
    27 => "01111", --   15
    28 => "01110", --   14
    29 => "01101", --   13
    30 => "01011", --   11
    31 => "01000", --    8
    32 => "00110", --    6
    33 => "00100", --    4
    34 => "00010", --    2
    35 => "11111", --   -1
    36 => "11101", --   -3
    37 => "11100", --   -4
    38 => "11010", --   -6
    39 => "11000", --   -8
    40 => "10111", --   -9
    41 => "10110", --  -10
    42 => "10101", --  -11
    43 => "10101", --  -11
    44 => "10100", --  -12
    45 => "10011", --  -13
    46 => "10011", --  -13
    47 => "10010", --  -14
    48 => "10001", --  -15
    49 => "10000", --  -16
    50 => "10000", --  -16
    51 => "10000", --  -16
    52 => "10000", --  -16
    53 => "10000", --  -16
    54 => "10000", --  -16
    55 => "10000", --  -16
    56 => "10000", --  -16
    57 => "10000", --  -16
    58 => "10000", --  -16
    59 => "10000", --  -16
    60 => "10000", --  -16
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  constant LUT_0_14_7_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11101", --   -3
    5 => "11101", --   -3
    6 => "11101", --   -3
    7 => "11101", --   -3
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11100", --   -4
    12 => "11011", --   -5
    13 => "11010", --   -6
    14 => "11010", --   -6
    15 => "11001", --   -7
    16 => "11000", --   -8
    17 => "11000", --   -8
    18 => "10111", --   -9
    19 => "10111", --   -9
    20 => "10111", --   -9
    21 => "10111", --   -9
    22 => "11000", --   -8
    23 => "11001", --   -7
    24 => "11010", --   -6
    25 => "11100", --   -4
    26 => "11101", --   -3
    27 => "11111", --   -1
    28 => "00000", --    0
    29 => "00010", --    2
    30 => "00011", --    3
    31 => "00100", --    4
    32 => "00101", --    5
    33 => "00110", --    6
    34 => "00110", --    6
    35 => "00110", --    6
    36 => "00110", --    6
    37 => "00110", --    6
    38 => "00101", --    5
    39 => "00100", --    4
    40 => "00011", --    3
    41 => "00011", --    3
    42 => "00010", --    2
    43 => "00001", --    1
    44 => "00000", --    0
    45 => "11111", --   -1
    46 => "11111", --   -1
    47 => "11110", --   -2
    48 => "11110", --   -2
    49 => "11110", --   -2
    50 => "11101", --   -3
    51 => "11101", --   -3
    52 => "11101", --   -3
    53 => "11101", --   -3
    54 => "11100", --   -4
    55 => "11100", --   -4
    56 => "11100", --   -4
    57 => "11011", --   -5
    58 => "11010", --   -6
    59 => "11001", --   -7
    60 => "11000", --   -8
    61 => "10111", --   -9
    62 => "10110", --  -10
    63 => "10101", --  -11
  );

  constant LUT_0_15_0_DATA : lut_array_t_0 := (
    0 => "11101", --   -3
    1 => "11101", --   -3
    2 => "11100", --   -4
    3 => "11011", --   -5
    4 => "11010", --   -6
    5 => "11001", --   -7
    6 => "11001", --   -7
    7 => "11000", --   -8
    8 => "10111", --   -9
    9 => "10111", --   -9
    10 => "10110", --  -10
    11 => "10110", --  -10
    12 => "10101", --  -11
    13 => "10101", --  -11
    14 => "10101", --  -11
    15 => "10101", --  -11
    16 => "10101", --  -11
    17 => "10110", --  -10
    18 => "10110", --  -10
    19 => "10111", --   -9
    20 => "11000", --   -8
    21 => "11001", --   -7
    22 => "11010", --   -6
    23 => "11011", --   -5
    24 => "11101", --   -3
    25 => "11110", --   -2
    26 => "11111", --   -1
    27 => "00000", --    0
    28 => "00001", --    1
    29 => "00001", --    1
    30 => "00010", --    2
    31 => "00011", --    3
    32 => "00011", --    3
    33 => "00011", --    3
    34 => "00100", --    4
    35 => "00100", --    4
    36 => "00100", --    4
    37 => "00100", --    4
    38 => "00100", --    4
    39 => "00101", --    5
    40 => "00101", --    5
    41 => "00101", --    5
    42 => "00110", --    6
    43 => "00110", --    6
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "01000", --    8
    47 => "01000", --    8
    48 => "01001", --    9
    49 => "01001", --    9
    50 => "01001", --    9
    51 => "01010", --   10
    52 => "01010", --   10
    53 => "01011", --   11
    54 => "01011", --   11
    55 => "01011", --   11
    56 => "01100", --   12
    57 => "01100", --   12
    58 => "01100", --   12
    59 => "01100", --   12
    60 => "01100", --   12
    61 => "01100", --   12
    62 => "01100", --   12
    63 => "01100", --   12
  );

  constant LUT_0_15_1_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11111", --   -1
    3 => "11111", --   -1
    4 => "11111", --   -1
    5 => "11111", --   -1
    6 => "11111", --   -1
    7 => "11111", --   -1
    8 => "11111", --   -1
    9 => "11111", --   -1
    10 => "11111", --   -1
    11 => "11111", --   -1
    12 => "11111", --   -1
    13 => "11111", --   -1
    14 => "11111", --   -1
    15 => "11110", --   -2
    16 => "11110", --   -2
    17 => "11110", --   -2
    18 => "11110", --   -2
    19 => "11110", --   -2
    20 => "11110", --   -2
    21 => "11110", --   -2
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11110", --   -2
    26 => "11111", --   -1
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "11111", --   -1
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "00000", --    0
    34 => "00001", --    1
    35 => "00001", --    1
    36 => "00001", --    1
    37 => "00010", --    2
    38 => "00010", --    2
    39 => "00011", --    3
    40 => "00011", --    3
    41 => "00011", --    3
    42 => "00100", --    4
    43 => "00100", --    4
    44 => "00101", --    5
    45 => "00101", --    5
    46 => "00110", --    6
    47 => "00110", --    6
    48 => "00111", --    7
    49 => "00111", --    7
    50 => "01000", --    8
    51 => "01000", --    8
    52 => "01001", --    9
    53 => "01001", --    9
    54 => "01010", --   10
    55 => "01010", --   10
    56 => "01011", --   11
    57 => "01100", --   12
    58 => "01100", --   12
    59 => "01101", --   13
    60 => "01101", --   13
    61 => "01110", --   14
    62 => "01110", --   14
    63 => "01111", --   15
  );

  constant LUT_0_15_2_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11101", --   -3
    3 => "11101", --   -3
    4 => "11100", --   -4
    5 => "11100", --   -4
    6 => "11011", --   -5
    7 => "11011", --   -5
    8 => "11010", --   -6
    9 => "11010", --   -6
    10 => "11010", --   -6
    11 => "11001", --   -7
    12 => "11001", --   -7
    13 => "11001", --   -7
    14 => "11001", --   -7
    15 => "11001", --   -7
    16 => "11010", --   -6
    17 => "11010", --   -6
    18 => "11010", --   -6
    19 => "11011", --   -5
    20 => "11011", --   -5
    21 => "11100", --   -4
    22 => "11100", --   -4
    23 => "11100", --   -4
    24 => "11101", --   -3
    25 => "11101", --   -3
    26 => "11110", --   -2
    27 => "11111", --   -1
    28 => "11111", --   -1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00001", --    1
    32 => "00010", --    2
    33 => "00010", --    2
    34 => "00011", --    3
    35 => "00011", --    3
    36 => "00100", --    4
    37 => "00100", --    4
    38 => "00101", --    5
    39 => "00101", --    5
    40 => "00110", --    6
    41 => "00110", --    6
    42 => "00110", --    6
    43 => "00111", --    7
    44 => "00111", --    7
    45 => "00111", --    7
    46 => "01000", --    8
    47 => "01000", --    8
    48 => "01000", --    8
    49 => "01000", --    8
    50 => "01001", --    9
    51 => "01001", --    9
    52 => "01001", --    9
    53 => "01010", --   10
    54 => "01010", --   10
    55 => "01011", --   11
    56 => "01011", --   11
    57 => "01100", --   12
    58 => "01100", --   12
    59 => "01101", --   13
    60 => "01101", --   13
    61 => "01110", --   14
    62 => "01110", --   14
    63 => "01110", --   14
  );

  constant LUT_0_15_3_DATA : lut_array_t_0 := (
    0 => "11100", --   -4
    1 => "11011", --   -5
    2 => "11010", --   -6
    3 => "11001", --   -7
    4 => "10111", --   -9
    5 => "10110", --  -10
    6 => "10101", --  -11
    7 => "10100", --  -12
    8 => "10011", --  -13
    9 => "10010", --  -14
    10 => "10010", --  -14
    11 => "10001", --  -15
    12 => "10001", --  -15
    13 => "10010", --  -14
    14 => "10010", --  -14
    15 => "10011", --  -13
    16 => "10011", --  -13
    17 => "10100", --  -12
    18 => "10101", --  -11
    19 => "10110", --  -10
    20 => "10111", --   -9
    21 => "11001", --   -7
    22 => "11010", --   -6
    23 => "11011", --   -5
    24 => "11100", --   -4
    25 => "11101", --   -3
    26 => "11101", --   -3
    27 => "11110", --   -2
    28 => "11111", --   -1
    29 => "00000", --    0
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00010", --    2
    33 => "00011", --    3
    34 => "00011", --    3
    35 => "00100", --    4
    36 => "00100", --    4
    37 => "00101", --    5
    38 => "00110", --    6
    39 => "00110", --    6
    40 => "00111", --    7
    41 => "01000", --    8
    42 => "01000", --    8
    43 => "01001", --    9
    44 => "01010", --   10
    45 => "01010", --   10
    46 => "01011", --   11
    47 => "01100", --   12
    48 => "01100", --   12
    49 => "01101", --   13
    50 => "01101", --   13
    51 => "01110", --   14
    52 => "01111", --   15
    53 => "01111", --   15
    54 => "01111", --   15
    55 => "01111", --   15
    56 => "01111", --   15
    57 => "01111", --   15
    58 => "01111", --   15
    59 => "01111", --   15
    60 => "01111", --   15
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_15_4_DATA : lut_array_t_0 := (
    0 => "11111", --   -1
    1 => "11111", --   -1
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11110", --   -2
    5 => "11110", --   -2
    6 => "11101", --   -3
    7 => "11101", --   -3
    8 => "11101", --   -3
    9 => "11100", --   -4
    10 => "11100", --   -4
    11 => "11100", --   -4
    12 => "11011", --   -5
    13 => "11011", --   -5
    14 => "11010", --   -6
    15 => "11010", --   -6
    16 => "11001", --   -7
    17 => "11001", --   -7
    18 => "11001", --   -7
    19 => "11000", --   -8
    20 => "11001", --   -7
    21 => "11001", --   -7
    22 => "11001", --   -7
    23 => "11010", --   -6
    24 => "11010", --   -6
    25 => "11011", --   -5
    26 => "11011", --   -5
    27 => "11100", --   -4
    28 => "11101", --   -3
    29 => "11110", --   -2
    30 => "11111", --   -1
    31 => "00000", --    0
    32 => "00001", --    1
    33 => "00001", --    1
    34 => "00010", --    2
    35 => "00011", --    3
    36 => "00100", --    4
    37 => "00101", --    5
    38 => "00110", --    6
    39 => "00111", --    7
    40 => "01000", --    8
    41 => "01001", --    9
    42 => "01001", --    9
    43 => "01010", --   10
    44 => "01011", --   11
    45 => "01100", --   12
    46 => "01100", --   12
    47 => "01101", --   13
    48 => "01101", --   13
    49 => "01110", --   14
    50 => "01110", --   14
    51 => "01111", --   15
    52 => "01111", --   15
    53 => "01111", --   15
    54 => "01111", --   15
    55 => "01110", --   14
    56 => "01110", --   14
    57 => "01110", --   14
    58 => "01110", --   14
    59 => "01110", --   14
    60 => "01110", --   14
    61 => "01111", --   15
    62 => "01111", --   15
    63 => "01111", --   15
  );

  constant LUT_0_15_5_DATA : lut_array_t_0 := (
    0 => "00001", --    1
    1 => "00010", --    2
    2 => "00010", --    2
    3 => "00010", --    2
    4 => "00011", --    3
    5 => "00011", --    3
    6 => "00011", --    3
    7 => "00011", --    3
    8 => "00011", --    3
    9 => "00100", --    4
    10 => "00100", --    4
    11 => "00100", --    4
    12 => "00100", --    4
    13 => "00100", --    4
    14 => "00100", --    4
    15 => "00100", --    4
    16 => "00011", --    3
    17 => "00011", --    3
    18 => "00011", --    3
    19 => "00011", --    3
    20 => "00010", --    2
    21 => "00010", --    2
    22 => "00010", --    2
    23 => "00010", --    2
    24 => "00001", --    1
    25 => "00001", --    1
    26 => "00001", --    1
    27 => "00001", --    1
    28 => "00001", --    1
    29 => "00000", --    0
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "00000", --    0
    33 => "11111", --   -1
    34 => "11111", --   -1
    35 => "11110", --   -2
    36 => "11110", --   -2
    37 => "11110", --   -2
    38 => "11101", --   -3
    39 => "11101", --   -3
    40 => "11101", --   -3
    41 => "11100", --   -4
    42 => "11100", --   -4
    43 => "11011", --   -5
    44 => "11011", --   -5
    45 => "11011", --   -5
    46 => "11010", --   -6
    47 => "11010", --   -6
    48 => "11010", --   -6
    49 => "11010", --   -6
    50 => "11001", --   -7
    51 => "11001", --   -7
    52 => "11001", --   -7
    53 => "11000", --   -8
    54 => "11000", --   -8
    55 => "11000", --   -8
    56 => "10111", --   -9
    57 => "10111", --   -9
    58 => "10110", --  -10
    59 => "10110", --  -10
    60 => "10110", --  -10
    61 => "10101", --  -11
    62 => "10101", --  -11
    63 => "10100", --  -12
  );

  constant LUT_0_15_6_DATA : lut_array_t_0 := (
    0 => "11110", --   -2
    1 => "11110", --   -2
    2 => "11110", --   -2
    3 => "11110", --   -2
    4 => "11101", --   -3
    5 => "11101", --   -3
    6 => "11101", --   -3
    7 => "11100", --   -4
    8 => "11100", --   -4
    9 => "11100", --   -4
    10 => "11011", --   -5
    11 => "11011", --   -5
    12 => "11011", --   -5
    13 => "11011", --   -5
    14 => "11011", --   -5
    15 => "11011", --   -5
    16 => "11011", --   -5
    17 => "11100", --   -4
    18 => "11100", --   -4
    19 => "11100", --   -4
    20 => "11101", --   -3
    21 => "11101", --   -3
    22 => "11110", --   -2
    23 => "11110", --   -2
    24 => "11110", --   -2
    25 => "11111", --   -1
    26 => "11111", --   -1
    27 => "00000", --    0
    28 => "00000", --    0
    29 => "00001", --    1
    30 => "00001", --    1
    31 => "00001", --    1
    32 => "00010", --    2
    33 => "00010", --    2
    34 => "00010", --    2
    35 => "00011", --    3
    36 => "00011", --    3
    37 => "00011", --    3
    38 => "00100", --    4
    39 => "00100", --    4
    40 => "00100", --    4
    41 => "00101", --    5
    42 => "00101", --    5
    43 => "00101", --    5
    44 => "00101", --    5
    45 => "00110", --    6
    46 => "00110", --    6
    47 => "00110", --    6
    48 => "00111", --    7
    49 => "00111", --    7
    50 => "00111", --    7
    51 => "01000", --    8
    52 => "01000", --    8
    53 => "01000", --    8
    54 => "01001", --    9
    55 => "01001", --    9
    56 => "01010", --   10
    57 => "01010", --   10
    58 => "01011", --   11
    59 => "01011", --   11
    60 => "01100", --   12
    61 => "01100", --   12
    62 => "01101", --   13
    63 => "01110", --   14
  );

  constant LUT_0_15_7_DATA : lut_array_t_0 := (
    0 => "00011", --    3
    1 => "00011", --    3
    2 => "00100", --    4
    3 => "00101", --    5
    4 => "00101", --    5
    5 => "00110", --    6
    6 => "00111", --    7
    7 => "00111", --    7
    8 => "01000", --    8
    9 => "01000", --    8
    10 => "01000", --    8
    11 => "01000", --    8
    12 => "01001", --    9
    13 => "01001", --    9
    14 => "01001", --    9
    15 => "01001", --    9
    16 => "01001", --    9
    17 => "01000", --    8
    18 => "01000", --    8
    19 => "01000", --    8
    20 => "00111", --    7
    21 => "00111", --    7
    22 => "00110", --    6
    23 => "00101", --    5
    24 => "00101", --    5
    25 => "00100", --    4
    26 => "00011", --    3
    27 => "00011", --    3
    28 => "00010", --    2
    29 => "00001", --    1
    30 => "00000", --    0
    31 => "00000", --    0
    32 => "11111", --   -1
    33 => "11110", --   -2
    34 => "11110", --   -2
    35 => "11101", --   -3
    36 => "11100", --   -4
    37 => "11100", --   -4
    38 => "11011", --   -5
    39 => "11011", --   -5
    40 => "11010", --   -6
    41 => "11001", --   -7
    42 => "11000", --   -8
    43 => "11000", --   -8
    44 => "10111", --   -9
    45 => "10111", --   -9
    46 => "10110", --  -10
    47 => "10101", --  -11
    48 => "10101", --  -11
    49 => "10100", --  -12
    50 => "10100", --  -12
    51 => "10011", --  -13
    52 => "10011", --  -13
    53 => "10011", --  -13
    54 => "10010", --  -14
    55 => "10010", --  -14
    56 => "10010", --  -14
    57 => "10001", --  -15
    58 => "10001", --  -15
    59 => "10001", --  -15
    60 => "10001", --  -15
    61 => "10000", --  -16
    62 => "10000", --  -16
    63 => "10000", --  -16
  );

  -- Layer 1 
  subtype  lut_array_t_1 is array (0 to 31) of signed(7 downto 0);

  constant LUT_1_0_0_DATA : lut_array_t_1 := (
    0 => "11010001", --  -47
    1 => "11010010", --  -46
    2 => "11010100", --  -44
    3 => "11010110", --  -42
    4 => "11011000", --  -40
    5 => "11011011", --  -37
    6 => "11011110", --  -34
    7 => "11100010", --  -30
    8 => "11100101", --  -27
    9 => "11100111", --  -25
    10 => "11101010", --  -22
    11 => "11101101", --  -19
    12 => "11101111", --  -17
    13 => "11110001", --  -15
    14 => "11110100", --  -12
    15 => "11110110", --  -10
    16 => "11111000", --   -8
    17 => "11111010", --   -6
    18 => "11111101", --   -3
    19 => "11111111", --   -1
    20 => "00000010", --    2
    21 => "00000100", --    4
    22 => "00000111", --    7
    23 => "00001010", --   10
    24 => "00001101", --   13
    25 => "00010001", --   17
    26 => "00010101", --   21
    27 => "00011001", --   25
    28 => "00011110", --   30
    29 => "00100010", --   34
    30 => "00100110", --   38
    31 => "00101010", --   42
  );

  constant LUT_1_0_1_DATA : lut_array_t_1 := (
    0 => "11011100", --  -36
    1 => "11011111", --  -33
    2 => "11100010", --  -30
    3 => "11100110", --  -26
    4 => "11101010", --  -22
    5 => "11101110", --  -18
    6 => "11110010", --  -14
    7 => "11110110", --  -10
    8 => "11111010", --   -6
    9 => "11111101", --   -3
    10 => "00000000", --    0
    11 => "00000010", --    2
    12 => "00000100", --    4
    13 => "00000110", --    6
    14 => "00001000", --    8
    15 => "00001001", --    9
    16 => "00001001", --    9
    17 => "00001010", --   10
    18 => "00001010", --   10
    19 => "00001001", --    9
    20 => "00001001", --    9
    21 => "00001000", --    8
    22 => "00000111", --    7
    23 => "00000110", --    6
    24 => "00000100", --    4
    25 => "00000011", --    3
    26 => "00000010", --    2
    27 => "00000001", --    1
    28 => "00000000", --    0
    29 => "11111111", --   -1
    30 => "11111101", --   -3
    31 => "11111101", --   -3
  );

  constant LUT_1_0_2_DATA : lut_array_t_1 := (
    0 => "00010111", --   23
    1 => "00010110", --   22
    2 => "00010101", --   21
    3 => "00010011", --   19
    4 => "00010010", --   18
    5 => "00010000", --   16
    6 => "00001110", --   14
    7 => "00001100", --   12
    8 => "00001010", --   10
    9 => "00001000", --    8
    10 => "00000110", --    6
    11 => "00000100", --    4
    12 => "00000001", --    1
    13 => "11111111", --   -1
    14 => "11111101", --   -3
    15 => "11111011", --   -5
    16 => "11111001", --   -7
    17 => "11111000", --   -8
    18 => "11110110", --  -10
    19 => "11110101", --  -11
    20 => "11110011", --  -13
    21 => "11110010", --  -14
    22 => "11110001", --  -15
    23 => "11101111", --  -17
    24 => "11101101", --  -19
    25 => "11101011", --  -21
    26 => "11101000", --  -24
    27 => "11100110", --  -26
    28 => "11100011", --  -29
    29 => "11100000", --  -32
    30 => "11011101", --  -35
    31 => "11011010", --  -38
  );

  constant LUT_1_0_3_DATA : lut_array_t_1 := (
    0 => "00000011", --    3
    1 => "00000100", --    4
    2 => "00000101", --    5
    3 => "00000101", --    5
    4 => "00000110", --    6
    5 => "00000110", --    6
    6 => "00000111", --    7
    7 => "00000111", --    7
    8 => "00000111", --    7
    9 => "00000111", --    7
    10 => "00000111", --    7
    11 => "00000111", --    7
    12 => "00000111", --    7
    13 => "00000111", --    7
    14 => "00000110", --    6
    15 => "00000110", --    6
    16 => "00000110", --    6
    17 => "00000101", --    5
    18 => "00000101", --    5
    19 => "00000100", --    4
    20 => "00000100", --    4
    21 => "00000011", --    3
    22 => "00000010", --    2
    23 => "00000001", --    1
    24 => "00000000", --    0
    25 => "11111110", --   -2
    26 => "11111101", --   -3
    27 => "11111011", --   -5
    28 => "11111001", --   -7
    29 => "11110111", --   -9
    30 => "11110101", --  -11
    31 => "11110011", --  -13
  );

  constant LUT_1_0_4_DATA : lut_array_t_1 := (
    0 => "11111100", --   -4
    1 => "11111011", --   -5
    2 => "11111011", --   -5
    3 => "11111011", --   -5
    4 => "11111011", --   -5
    5 => "11111011", --   -5
    6 => "11111011", --   -5
    7 => "11111011", --   -5
    8 => "11111100", --   -4
    9 => "11111100", --   -4
    10 => "11111100", --   -4
    11 => "11111101", --   -3
    12 => "11111101", --   -3
    13 => "11111110", --   -2
    14 => "11111111", --   -1
    15 => "11111111", --   -1
    16 => "00000000", --    0
    17 => "00000000", --    0
    18 => "00000001", --    1
    19 => "00000001", --    1
    20 => "00000010", --    2
    21 => "00000010", --    2
    22 => "00000010", --    2
    23 => "00000010", --    2
    24 => "00000010", --    2
    25 => "00000010", --    2
    26 => "00000010", --    2
    27 => "00000010", --    2
    28 => "00000010", --    2
    29 => "00000010", --    2
    30 => "00000010", --    2
    31 => "00000010", --    2
  );

  constant LUT_1_1_0_DATA : lut_array_t_1 := (
    0 => "11110110", --  -10
    1 => "11110110", --  -10
    2 => "11110110", --  -10
    3 => "11110110", --  -10
    4 => "11110101", --  -11
    5 => "11110101", --  -11
    6 => "11110101", --  -11
    7 => "11110110", --  -10
    8 => "11110110", --  -10
    9 => "11110110", --  -10
    10 => "11110111", --   -9
    11 => "11110111", --   -9
    12 => "11111000", --   -8
    13 => "11111001", --   -7
    14 => "11111010", --   -6
    15 => "11111011", --   -5
    16 => "11111100", --   -4
    17 => "11111101", --   -3
    18 => "11111110", --   -2
    19 => "00000000", --    0
    20 => "00000001", --    1
    21 => "00000011", --    3
    22 => "00000100", --    4
    23 => "00000110", --    6
    24 => "00001000", --    8
    25 => "00001001", --    9
    26 => "00001011", --   11
    27 => "00001101", --   13
    28 => "00001110", --   14
    29 => "00010000", --   16
    30 => "00010001", --   17
    31 => "00010011", --   19
  );

  constant LUT_1_1_1_DATA : lut_array_t_1 := (
    0 => "00000100", --    4
    1 => "00000100", --    4
    2 => "00000011", --    3
    3 => "00000011", --    3
    4 => "00000011", --    3
    5 => "00000010", --    2
    6 => "00000010", --    2
    7 => "00000001", --    1
    8 => "00000001", --    1
    9 => "00000000", --    0
    10 => "11111111", --   -1
    11 => "11111111", --   -1
    12 => "11111110", --   -2
    13 => "11111110", --   -2
    14 => "11111110", --   -2
    15 => "11111110", --   -2
    16 => "11111110", --   -2
    17 => "11111110", --   -2
    18 => "11111111", --   -1
    19 => "11111111", --   -1
    20 => "00000000", --    0
    21 => "00000001", --    1
    22 => "00000001", --    1
    23 => "00000010", --    2
    24 => "00000011", --    3
    25 => "00000011", --    3
    26 => "00000011", --    3
    27 => "00000100", --    4
    28 => "00000100", --    4
    29 => "00000100", --    4
    30 => "00000100", --    4
    31 => "00000011", --    3
  );

  constant LUT_1_1_2_DATA : lut_array_t_1 := (
    0 => "11010010", --  -46
    1 => "11010010", --  -46
    2 => "11010100", --  -44
    3 => "11010110", --  -42
    4 => "11011001", --  -39
    5 => "11011101", --  -35
    6 => "11100001", --  -31
    7 => "11100101", --  -27
    8 => "11101010", --  -22
    9 => "11101111", --  -17
    10 => "11110100", --  -12
    11 => "11111000", --   -8
    12 => "11111101", --   -3
    13 => "00000001", --    1
    14 => "00000101", --    5
    15 => "00001000", --    8
    16 => "00001010", --   10
    17 => "00001011", --   11
    18 => "00001100", --   12
    19 => "00001100", --   12
    20 => "00001011", --   11
    21 => "00001001", --    9
    22 => "00000111", --    7
    23 => "00000101", --    5
    24 => "00000010", --    2
    25 => "11111111", --   -1
    26 => "11111100", --   -4
    27 => "11111001", --   -7
    28 => "11110110", --  -10
    29 => "11110011", --  -13
    30 => "11110001", --  -15
    31 => "11101111", --  -17
  );

  constant LUT_1_1_3_DATA : lut_array_t_1 := (
    0 => "11111000", --   -8
    1 => "11111011", --   -5
    2 => "11111101", --   -3
    3 => "00000000", --    0
    4 => "00000011", --    3
    5 => "00000101", --    5
    6 => "00001000", --    8
    7 => "00001001", --    9
    8 => "00001011", --   11
    9 => "00001011", --   11
    10 => "00001011", --   11
    11 => "00001011", --   11
    12 => "00001011", --   11
    13 => "00001010", --   10
    14 => "00001001", --    9
    15 => "00001000", --    8
    16 => "00000110", --    6
    17 => "00000101", --    5
    18 => "00000011", --    3
    19 => "00000010", --    2
    20 => "00000000", --    0
    21 => "11111111", --   -1
    22 => "11111101", --   -3
    23 => "11111100", --   -4
    24 => "11111010", --   -6
    25 => "11111001", --   -7
    26 => "11110111", --   -9
    27 => "11110110", --  -10
    28 => "11110101", --  -11
    29 => "11110100", --  -12
    30 => "11110011", --  -13
    31 => "11110010", --  -14
  );

  constant LUT_1_1_4_DATA : lut_array_t_1 := (
    0 => "00010001", --   17
    1 => "00010000", --   16
    2 => "00010000", --   16
    3 => "00001111", --   15
    4 => "00001110", --   14
    5 => "00001101", --   13
    6 => "00001100", --   12
    7 => "00001010", --   10
    8 => "00001001", --    9
    9 => "00000111", --    7
    10 => "00000101", --    5
    11 => "00000011", --    3
    12 => "00000001", --    1
    13 => "11111110", --   -2
    14 => "11111100", --   -4
    15 => "11111010", --   -6
    16 => "11111000", --   -8
    17 => "11110111", --   -9
    18 => "11110101", --  -11
    19 => "11110011", --  -13
    20 => "11110010", --  -14
    21 => "11110001", --  -15
    22 => "11110000", --  -16
    23 => "11101111", --  -17
    24 => "11101110", --  -18
    25 => "11101110", --  -18
    26 => "11101110", --  -18
    27 => "11101101", --  -19
    28 => "11101101", --  -19
    29 => "11101110", --  -18
    30 => "11101110", --  -18
    31 => "11101110", --  -18
  );

  constant LUT_1_2_0_DATA : lut_array_t_1 := (
    0 => "11100100", --  -28
    1 => "11100101", --  -27
    2 => "11100110", --  -26
    3 => "11100111", --  -25
    4 => "11100111", --  -25
    5 => "11101000", --  -24
    6 => "11101001", --  -23
    7 => "11101010", --  -22
    8 => "11101010", --  -22
    9 => "11101011", --  -21
    10 => "11101011", --  -21
    11 => "11101100", --  -20
    12 => "11101101", --  -19
    13 => "11101110", --  -18
    14 => "11101111", --  -17
    15 => "11110000", --  -16
    16 => "11110010", --  -14
    17 => "11110101", --  -11
    18 => "11111000", --   -8
    19 => "11111011", --   -5
    20 => "11111111", --   -1
    21 => "00000011", --    3
    22 => "00001000", --    8
    23 => "00001101", --   13
    24 => "00010010", --   18
    25 => "00011000", --   24
    26 => "00011111", --   31
    27 => "00100101", --   37
    28 => "00101100", --   44
    29 => "00110011", --   51
    30 => "00111001", --   57
    31 => "01000000", --   64
  );

  constant LUT_1_2_1_DATA : lut_array_t_1 := (
    0 => "00011011", --   27
    1 => "00011010", --   26
    2 => "00011001", --   25
    3 => "00011000", --   24
    4 => "00010111", --   23
    5 => "00010101", --   21
    6 => "00010011", --   19
    7 => "00010001", --   17
    8 => "00001111", --   15
    9 => "00001100", --   12
    10 => "00001010", --   10
    11 => "00000111", --    7
    12 => "00000100", --    4
    13 => "00000010", --    2
    14 => "11111111", --   -1
    15 => "11111101", --   -3
    16 => "11111011", --   -5
    17 => "11111001", --   -7
    18 => "11110111", --   -9
    19 => "11110110", --  -10
    20 => "11110100", --  -12
    21 => "11110011", --  -13
    22 => "11110010", --  -14
    23 => "11110000", --  -16
    24 => "11101111", --  -17
    25 => "11101101", --  -19
    26 => "11101100", --  -20
    27 => "11101010", --  -22
    28 => "11101000", --  -24
    29 => "11100110", --  -26
    30 => "11100011", --  -29
    31 => "11100001", --  -31
  );

  constant LUT_1_2_2_DATA : lut_array_t_1 := (
    0 => "11110101", --  -11
    1 => "11110110", --  -10
    2 => "11110111", --   -9
    3 => "11111000", --   -8
    4 => "11111010", --   -6
    5 => "11111011", --   -5
    6 => "11111100", --   -4
    7 => "11111110", --   -2
    8 => "11111111", --   -1
    9 => "00000001", --    1
    10 => "00000010", --    2
    11 => "00000100", --    4
    12 => "00000101", --    5
    13 => "00000110", --    6
    14 => "00000111", --    7
    15 => "00000111", --    7
    16 => "00000111", --    7
    17 => "00000111", --    7
    18 => "00000110", --    6
    19 => "00000100", --    4
    20 => "00000011", --    3
    21 => "00000001", --    1
    22 => "11111110", --   -2
    23 => "11111011", --   -5
    24 => "11111000", --   -8
    25 => "11110100", --  -12
    26 => "11110000", --  -16
    27 => "11101100", --  -20
    28 => "11101000", --  -24
    29 => "11100011", --  -29
    30 => "11100000", --  -32
    31 => "11011100", --  -36
  );

  constant LUT_1_2_3_DATA : lut_array_t_1 := (
    0 => "11111001", --   -7
    1 => "11111001", --   -7
    2 => "11111010", --   -6
    3 => "11111011", --   -5
    4 => "11111100", --   -4
    5 => "11111101", --   -3
    6 => "11111110", --   -2
    7 => "00000000", --    0
    8 => "00000001", --    1
    9 => "00000010", --    2
    10 => "00000011", --    3
    11 => "00000100", --    4
    12 => "00000110", --    6
    13 => "00000111", --    7
    14 => "00001000", --    8
    15 => "00001001", --    9
    16 => "00001010", --   10
    17 => "00001010", --   10
    18 => "00001011", --   11
    19 => "00001011", --   11
    20 => "00001010", --   10
    21 => "00001010", --   10
    22 => "00001000", --    8
    23 => "00000110", --    6
    24 => "00000011", --    3
    25 => "00000000", --    0
    26 => "11111011", --   -5
    27 => "11110110", --  -10
    28 => "11110001", --  -15
    29 => "11101011", --  -21
    30 => "11100110", --  -26
    31 => "11100001", --  -31
  );

  constant LUT_1_2_4_DATA : lut_array_t_1 := (
    0 => "00000101", --    5
    1 => "00000110", --    6
    2 => "00000111", --    7
    3 => "00000111", --    7
    4 => "00001000", --    8
    5 => "00001000", --    8
    6 => "00001000", --    8
    7 => "00001000", --    8
    8 => "00001000", --    8
    9 => "00000111", --    7
    10 => "00000111", --    7
    11 => "00000110", --    6
    12 => "00000101", --    5
    13 => "00000100", --    4
    14 => "00000011", --    3
    15 => "00000010", --    2
    16 => "00000001", --    1
    17 => "00000000", --    0
    18 => "11111111", --   -1
    19 => "11111110", --   -2
    20 => "11111101", --   -3
    21 => "11111100", --   -4
    22 => "11111100", --   -4
    23 => "11111011", --   -5
    24 => "11111010", --   -6
    25 => "11111010", --   -6
    26 => "11111001", --   -7
    27 => "11111000", --   -8
    28 => "11111000", --   -8
    29 => "11110111", --   -9
    30 => "11110110", --  -10
    31 => "11110110", --  -10
  );

  constant LUT_1_3_0_DATA : lut_array_t_1 := (
    0 => "11100111", --  -25
    1 => "11101001", --  -23
    2 => "11101011", --  -21
    3 => "11101101", --  -19
    4 => "11101111", --  -17
    5 => "11110010", --  -14
    6 => "11110100", --  -12
    7 => "11110111", --   -9
    8 => "11111001", --   -7
    9 => "11111011", --   -5
    10 => "11111101", --   -3
    11 => "11111111", --   -1
    12 => "00000001", --    1
    13 => "00000010", --    2
    14 => "00000011", --    3
    15 => "00000100", --    4
    16 => "00000101", --    5
    17 => "00000110", --    6
    18 => "00000110", --    6
    19 => "00000110", --    6
    20 => "00000110", --    6
    21 => "00000110", --    6
    22 => "00000110", --    6
    23 => "00000110", --    6
    24 => "00000110", --    6
    25 => "00000110", --    6
    26 => "00000110", --    6
    27 => "00000110", --    6
    28 => "00000110", --    6
    29 => "00000110", --    6
    30 => "00000111", --    7
    31 => "00000111", --    7
  );

  constant LUT_1_3_1_DATA : lut_array_t_1 := (
    0 => "00010001", --   17
    1 => "00010000", --   16
    2 => "00001111", --   15
    3 => "00001101", --   13
    4 => "00001100", --   12
    5 => "00001011", --   11
    6 => "00001001", --    9
    7 => "00001000", --    8
    8 => "00000110", --    6
    9 => "00000101", --    5
    10 => "00000100", --    4
    11 => "00000010", --    2
    12 => "00000001", --    1
    13 => "00000000", --    0
    14 => "11111111", --   -1
    15 => "11111110", --   -2
    16 => "11111100", --   -4
    17 => "11111011", --   -5
    18 => "11111010", --   -6
    19 => "11111001", --   -7
    20 => "11111000", --   -8
    21 => "11111000", --   -8
    22 => "11110111", --   -9
    23 => "11110110", --  -10
    24 => "11110101", --  -11
    25 => "11110100", --  -12
    26 => "11110011", --  -13
    27 => "11110010", --  -14
    28 => "11110000", --  -16
    29 => "11110000", --  -16
    30 => "11101111", --  -17
    31 => "11101110", --  -18
  );

  constant LUT_1_3_2_DATA : lut_array_t_1 := (
    0 => "11111111", --   -1
    1 => "00000000", --    0
    2 => "00000001", --    1
    3 => "00000010", --    2
    4 => "00000011", --    3
    5 => "00000100", --    4
    6 => "00000101", --    5
    7 => "00000110", --    6
    8 => "00000110", --    6
    9 => "00000111", --    7
    10 => "00000111", --    7
    11 => "00000111", --    7
    12 => "00000110", --    6
    13 => "00000110", --    6
    14 => "00000101", --    5
    15 => "00000100", --    4
    16 => "00000011", --    3
    17 => "00000010", --    2
    18 => "00000001", --    1
    19 => "11111111", --   -1
    20 => "11111101", --   -3
    21 => "11111011", --   -5
    22 => "11111010", --   -6
    23 => "11111000", --   -8
    24 => "11110110", --  -10
    25 => "11110100", --  -12
    26 => "11110010", --  -14
    27 => "11110001", --  -15
    28 => "11101111", --  -17
    29 => "11101110", --  -18
    30 => "11101101", --  -19
    31 => "11101100", --  -20
  );

  constant LUT_1_3_3_DATA : lut_array_t_1 := (
    0 => "00010010", --   18
    1 => "00010001", --   17
    2 => "00010001", --   17
    3 => "00010001", --   17
    4 => "00010001", --   17
    5 => "00010000", --   16
    6 => "00010000", --   16
    7 => "00001111", --   15
    8 => "00001110", --   14
    9 => "00001101", --   13
    10 => "00001100", --   12
    11 => "00001011", --   11
    12 => "00001010", --   10
    13 => "00001000", --    8
    14 => "00000110", --    6
    15 => "00000100", --    4
    16 => "00000010", --    2
    17 => "00000000", --    0
    18 => "11111110", --   -2
    19 => "11111011", --   -5
    20 => "11111001", --   -7
    21 => "11110110", --  -10
    22 => "11110100", --  -12
    23 => "11110001", --  -15
    24 => "11101111", --  -17
    25 => "11101101", --  -19
    26 => "11101011", --  -21
    27 => "11101001", --  -23
    28 => "11100111", --  -25
    29 => "11100101", --  -27
    30 => "11100011", --  -29
    31 => "11100010", --  -30
  );

  constant LUT_1_3_4_DATA : lut_array_t_1 := (
    0 => "11000000", --  -64
    1 => "11000001", --  -63
    2 => "11000010", --  -62
    3 => "11000100", --  -60
    4 => "11000111", --  -57
    5 => "11001010", --  -54
    6 => "11001101", --  -51
    7 => "11010001", --  -47
    8 => "11010101", --  -43
    9 => "11011001", --  -39
    10 => "11011101", --  -35
    11 => "11100010", --  -30
    12 => "11100110", --  -26
    13 => "11101010", --  -22
    14 => "11101111", --  -17
    15 => "11110011", --  -13
    16 => "11110111", --   -9
    17 => "11111011", --   -5
    18 => "00000000", --    0
    19 => "00000100", --    4
    20 => "00001000", --    8
    21 => "00001011", --   11
    22 => "00001111", --   15
    23 => "00010011", --   19
    24 => "00010110", --   22
    25 => "00011001", --   25
    26 => "00011100", --   28
    27 => "00011111", --   31
    28 => "00100001", --   33
    29 => "00100100", --   36
    30 => "00100110", --   38
    31 => "00101000", --   40
  );

  constant LUT_1_4_0_DATA : lut_array_t_1 := (
    0 => "11100010", --  -30
    1 => "11100001", --  -31
    2 => "11100000", --  -32
    3 => "11100000", --  -32
    4 => "11100000", --  -32
    5 => "11100001", --  -31
    6 => "11100001", --  -31
    7 => "11100010", --  -30
    8 => "11100100", --  -28
    9 => "11100101", --  -27
    10 => "11100111", --  -25
    11 => "11101001", --  -23
    12 => "11101011", --  -21
    13 => "11101110", --  -18
    14 => "11110000", --  -16
    15 => "11110011", --  -13
    16 => "11110101", --  -11
    17 => "11111000", --   -8
    18 => "11111011", --   -5
    19 => "11111101", --   -3
    20 => "00000000", --    0
    21 => "00000010", --    2
    22 => "00000101", --    5
    23 => "00000111", --    7
    24 => "00001001", --    9
    25 => "00001010", --   10
    26 => "00001100", --   12
    27 => "00001101", --   13
    28 => "00001110", --   14
    29 => "00001111", --   15
    30 => "00010000", --   16
    31 => "00010000", --   16
  );

  constant LUT_1_4_1_DATA : lut_array_t_1 := (
    0 => "11110001", --  -15
    1 => "11110001", --  -15
    2 => "11110010", --  -14
    3 => "11110011", --  -13
    4 => "11110100", --  -12
    5 => "11110101", --  -11
    6 => "11110111", --   -9
    7 => "11111000", --   -8
    8 => "11111010", --   -6
    9 => "11111011", --   -5
    10 => "11111101", --   -3
    11 => "11111110", --   -2
    12 => "11111111", --   -1
    13 => "00000000", --    0
    14 => "00000001", --    1
    15 => "00000010", --    2
    16 => "00000010", --    2
    17 => "00000010", --    2
    18 => "00000010", --    2
    19 => "00000001", --    1
    20 => "00000000", --    0
    21 => "00000000", --    0
    22 => "11111111", --   -1
    23 => "11111110", --   -2
    24 => "11111101", --   -3
    25 => "11111100", --   -4
    26 => "11111011", --   -5
    27 => "11111011", --   -5
    28 => "11111010", --   -6
    29 => "11111001", --   -7
    30 => "11111001", --   -7
    31 => "11111000", --   -8
  );

  constant LUT_1_4_2_DATA : lut_array_t_1 := (
    0 => "00001011", --   11
    1 => "00001011", --   11
    2 => "00001100", --   12
    3 => "00001101", --   13
    4 => "00001110", --   14
    5 => "00001110", --   14
    6 => "00001110", --   14
    7 => "00001110", --   14
    8 => "00001110", --   14
    9 => "00001101", --   13
    10 => "00001100", --   12
    11 => "00001011", --   11
    12 => "00001001", --    9
    13 => "00000111", --    7
    14 => "00000101", --    5
    15 => "00000011", --    3
    16 => "00000000", --    0
    17 => "11111110", --   -2
    18 => "11111011", --   -5
    19 => "11111000", --   -8
    20 => "11110101", --  -11
    21 => "11110010", --  -14
    22 => "11101111", --  -17
    23 => "11101101", --  -19
    24 => "11101010", --  -22
    25 => "11101000", --  -24
    26 => "11100110", --  -26
    27 => "11100101", --  -27
    28 => "11100100", --  -28
    29 => "11100011", --  -29
    30 => "11100010", --  -30
    31 => "11100001", --  -31
  );

  constant LUT_1_4_3_DATA : lut_array_t_1 := (
    0 => "00100011", --   35
    1 => "00100010", --   34
    2 => "00100001", --   33
    3 => "00011111", --   31
    4 => "00011110", --   30
    5 => "00011100", --   28
    6 => "00011001", --   25
    7 => "00010111", --   23
    8 => "00010100", --   20
    9 => "00010010", --   18
    10 => "00001111", --   15
    11 => "00001100", --   12
    12 => "00001001", --    9
    13 => "00000110", --    6
    14 => "00000011", --    3
    15 => "00000000", --    0
    16 => "11111101", --   -3
    17 => "11111010", --   -6
    18 => "11111000", --   -8
    19 => "11110101", --  -11
    20 => "11110010", --  -14
    21 => "11110000", --  -16
    22 => "11101101", --  -19
    23 => "11101010", --  -22
    24 => "11100111", --  -25
    25 => "11100100", --  -28
    26 => "11100001", --  -31
    27 => "11011101", --  -35
    28 => "11011010", --  -38
    29 => "11010110", --  -42
    30 => "11010011", --  -45
    31 => "11001111", --  -49
  );

  constant LUT_1_4_4_DATA : lut_array_t_1 := (
    0 => "11011100", --  -36
    1 => "11011101", --  -35
    2 => "11100000", --  -32
    3 => "11100011", --  -29
    4 => "11100111", --  -25
    5 => "11101010", --  -22
    6 => "11101110", --  -18
    7 => "11110011", --  -13
    8 => "11110110", --  -10
    9 => "11111010", --   -6
    10 => "11111101", --   -3
    11 => "00000000", --    0
    12 => "00000011", --    3
    13 => "00000101", --    5
    14 => "00000111", --    7
    15 => "00001000", --    8
    16 => "00001001", --    9
    17 => "00001010", --   10
    18 => "00001001", --    9
    19 => "00001001", --    9
    20 => "00001000", --    8
    21 => "00000111", --    7
    22 => "00000101", --    5
    23 => "00000011", --    3
    24 => "00000010", --    2
    25 => "00000000", --    0
    26 => "11111110", --   -2
    27 => "11111100", --   -4
    28 => "11111011", --   -5
    29 => "11111001", --   -7
    30 => "11110111", --   -9
    31 => "11110101", --  -11
  );

  constant LUT_1_5_0_DATA : lut_array_t_1 := (
    0 => "00001001", --    9
    1 => "00001001", --    9
    2 => "00001010", --   10
    3 => "00001011", --   11
    4 => "00001011", --   11
    5 => "00001100", --   12
    6 => "00001100", --   12
    7 => "00001100", --   12
    8 => "00001100", --   12
    9 => "00001100", --   12
    10 => "00001011", --   11
    11 => "00001010", --   10
    12 => "00001001", --    9
    13 => "00001000", --    8
    14 => "00000111", --    7
    15 => "00000101", --    5
    16 => "00000100", --    4
    17 => "00000010", --    2
    18 => "00000001", --    1
    19 => "11111111", --   -1
    20 => "11111101", --   -3
    21 => "11111100", --   -4
    22 => "11111010", --   -6
    23 => "11111001", --   -7
    24 => "11110111", --   -9
    25 => "11110110", --  -10
    26 => "11110101", --  -11
    27 => "11110011", --  -13
    28 => "11110010", --  -14
    29 => "11110001", --  -15
    30 => "11110000", --  -16
    31 => "11101111", --  -17
  );

  constant LUT_1_5_1_DATA : lut_array_t_1 := (
    0 => "00001111", --   15
    1 => "00001110", --   14
    2 => "00001101", --   13
    3 => "00001100", --   12
    4 => "00001010", --   10
    5 => "00001001", --    9
    6 => "00001000", --    8
    7 => "00000110", --    6
    8 => "00000101", --    5
    9 => "00000011", --    3
    10 => "00000010", --    2
    11 => "00000000", --    0
    12 => "11111111", --   -1
    13 => "11111101", --   -3
    14 => "11111100", --   -4
    15 => "11111100", --   -4
    16 => "11111011", --   -5
    17 => "11111011", --   -5
    18 => "11111011", --   -5
    19 => "11111011", --   -5
    20 => "11111100", --   -4
    21 => "11111101", --   -3
    22 => "11111101", --   -3
    23 => "11111110", --   -2
    24 => "11111111", --   -1
    25 => "00000000", --    0
    26 => "00000001", --    1
    27 => "00000010", --    2
    28 => "00000011", --    3
    29 => "00000100", --    4
    30 => "00000101", --    5
    31 => "00000110", --    6
  );

  constant LUT_1_5_2_DATA : lut_array_t_1 := (
    0 => "11000001", --  -63
    1 => "11000001", --  -63
    2 => "11000010", --  -62
    3 => "11000100", --  -60
    4 => "11000110", --  -58
    5 => "11001001", --  -55
    6 => "11001101", --  -51
    7 => "11010001", --  -47
    8 => "11010110", --  -42
    9 => "11011100", --  -36
    10 => "11100001", --  -31
    11 => "11101000", --  -24
    12 => "11101110", --  -18
    13 => "11110100", --  -12
    14 => "11111010", --   -6
    15 => "00000000", --    0
    16 => "00000110", --    6
    17 => "00001011", --   11
    18 => "00010000", --   16
    19 => "00010100", --   20
    20 => "00011000", --   24
    21 => "00011011", --   27
    22 => "00011101", --   29
    23 => "00011111", --   31
    24 => "00011111", --   31
    25 => "00100000", --   32
    26 => "00011111", --   31
    27 => "00011110", --   30
    28 => "00011100", --   28
    29 => "00011010", --   26
    30 => "00011001", --   25
    31 => "00010111", --   23
  );

  constant LUT_1_5_3_DATA : lut_array_t_1 := (
    0 => "11110011", --  -13
    1 => "11111001", --   -7
    2 => "11111111", --   -1
    3 => "00000101", --    5
    4 => "00001010", --   10
    5 => "00001111", --   15
    6 => "00010011", --   19
    7 => "00010110", --   22
    8 => "00011000", --   24
    9 => "00011001", --   25
    10 => "00011001", --   25
    11 => "00011000", --   24
    12 => "00010110", --   22
    13 => "00010100", --   20
    14 => "00010001", --   17
    15 => "00001110", --   14
    16 => "00001010", --   10
    17 => "00000110", --    6
    18 => "00000001", --    1
    19 => "11111101", --   -3
    20 => "11111001", --   -7
    21 => "11110101", --  -11
    22 => "11110001", --  -15
    23 => "11101110", --  -18
    24 => "11101100", --  -20
    25 => "11101010", --  -22
    26 => "11101010", --  -22
    27 => "11101010", --  -22
    28 => "11101010", --  -22
    29 => "11101011", --  -21
    30 => "11101100", --  -20
    31 => "11101101", --  -19
  );

  constant LUT_1_5_4_DATA : lut_array_t_1 := (
    0 => "00000101", --    5
    1 => "00000100", --    4
    2 => "00000011", --    3
    3 => "00000010", --    2
    4 => "00000001", --    1
    5 => "00000000", --    0
    6 => "11111111", --   -1
    7 => "11111110", --   -2
    8 => "11111110", --   -2
    9 => "11111101", --   -3
    10 => "11111101", --   -3
    11 => "11111101", --   -3
    12 => "11111101", --   -3
    13 => "11111101", --   -3
    14 => "11111101", --   -3
    15 => "11111101", --   -3
    16 => "11111101", --   -3
    17 => "11111101", --   -3
    18 => "11111101", --   -3
    19 => "11111110", --   -2
    20 => "11111110", --   -2
    21 => "11111110", --   -2
    22 => "11111110", --   -2
    23 => "11111110", --   -2
    24 => "11111111", --   -1
    25 => "11111111", --   -1
    26 => "11111111", --   -1
    27 => "11111111", --   -1
    28 => "11111111", --   -1
    29 => "11111111", --   -1
    30 => "11111110", --   -2
    31 => "11111110", --   -2
  );

  constant LUT_1_6_0_DATA : lut_array_t_1 := (
    0 => "00001000", --    8
    1 => "00001000", --    8
    2 => "00001001", --    9
    3 => "00001001", --    9
    4 => "00001001", --    9
    5 => "00001001", --    9
    6 => "00001001", --    9
    7 => "00001000", --    8
    8 => "00000111", --    7
    9 => "00000110", --    6
    10 => "00000100", --    4
    11 => "00000010", --    2
    12 => "00000000", --    0
    13 => "11111110", --   -2
    14 => "11111100", --   -4
    15 => "11111010", --   -6
    16 => "11111000", --   -8
    17 => "11110110", --  -10
    18 => "11110101", --  -11
    19 => "11110100", --  -12
    20 => "11110010", --  -14
    21 => "11110010", --  -14
    22 => "11110001", --  -15
    23 => "11110001", --  -15
    24 => "11110001", --  -15
    25 => "11110001", --  -15
    26 => "11110010", --  -14
    27 => "11110010", --  -14
    28 => "11110011", --  -13
    29 => "11110100", --  -12
    30 => "11110101", --  -11
    31 => "11110110", --  -10
  );

  constant LUT_1_6_1_DATA : lut_array_t_1 := (
    0 => "00000010", --    2
    1 => "00000001", --    1
    2 => "00000001", --    1
    3 => "00000000", --    0
    4 => "11111111", --   -1
    5 => "11111110", --   -2
    6 => "11111101", --   -3
    7 => "11111100", --   -4
    8 => "11111011", --   -5
    9 => "11111001", --   -7
    10 => "11111000", --   -8
    11 => "11110110", --  -10
    12 => "11110101", --  -11
    13 => "11110100", --  -12
    14 => "11110100", --  -12
    15 => "11110100", --  -12
    16 => "11110101", --  -11
    17 => "11110110", --  -10
    18 => "11111000", --   -8
    19 => "11111010", --   -6
    20 => "11111101", --   -3
    21 => "00000000", --    0
    22 => "00000011", --    3
    23 => "00000110", --    6
    24 => "00001001", --    9
    25 => "00001011", --   11
    26 => "00001110", --   14
    27 => "00010000", --   16
    28 => "00010010", --   18
    29 => "00010011", --   19
    30 => "00010101", --   21
    31 => "00010110", --   22
  );

  constant LUT_1_6_2_DATA : lut_array_t_1 := (
    0 => "11111010", --   -6
    1 => "11111010", --   -6
    2 => "11111010", --   -6
    3 => "11111010", --   -6
    4 => "11111011", --   -5
    5 => "11111100", --   -4
    6 => "11111101", --   -3
    7 => "11111110", --   -2
    8 => "00000000", --    0
    9 => "00000010", --    2
    10 => "00000100", --    4
    11 => "00000110", --    6
    12 => "00001000", --    8
    13 => "00001001", --    9
    14 => "00001010", --   10
    15 => "00001010", --   10
    16 => "00001001", --    9
    17 => "00001000", --    8
    18 => "00000101", --    5
    19 => "00000010", --    2
    20 => "11111110", --   -2
    21 => "11111001", --   -7
    22 => "11110100", --  -12
    23 => "11101111", --  -17
    24 => "11101001", --  -23
    25 => "11100100", --  -28
    26 => "11011110", --  -34
    27 => "11011001", --  -39
    28 => "11010100", --  -44
    29 => "11010000", --  -48
    30 => "11001100", --  -52
    31 => "11001000", --  -56
  );

  constant LUT_1_6_3_DATA : lut_array_t_1 := (
    0 => "00000011", --    3
    1 => "00000011", --    3
    2 => "00000011", --    3
    3 => "00000011", --    3
    4 => "00000011", --    3
    5 => "00000011", --    3
    6 => "00000011", --    3
    7 => "00000100", --    4
    8 => "00000100", --    4
    9 => "00000101", --    5
    10 => "00000110", --    6
    11 => "00000111", --    7
    12 => "00001000", --    8
    13 => "00001001", --    9
    14 => "00001010", --   10
    15 => "00001011", --   11
    16 => "00001100", --   12
    17 => "00001100", --   12
    18 => "00001101", --   13
    19 => "00001100", --   12
    20 => "00001100", --   12
    21 => "00001010", --   10
    22 => "00001000", --    8
    23 => "00000101", --    5
    24 => "00000000", --    0
    25 => "11111010", --   -6
    26 => "11110100", --  -12
    27 => "11101100", --  -20
    28 => "11100011", --  -29
    29 => "11011011", --  -37
    30 => "11010010", --  -46
    31 => "11001001", --  -55
  );

  constant LUT_1_6_4_DATA : lut_array_t_1 := (
    0 => "11011111", --  -33
    1 => "11011111", --  -33
    2 => "11011111", --  -33
    3 => "11011111", --  -33
    4 => "11011111", --  -33
    5 => "11011111", --  -33
    6 => "11011111", --  -33
    7 => "11011111", --  -33
    8 => "11011111", --  -33
    9 => "11011111", --  -33
    10 => "11011111", --  -33
    11 => "11011111", --  -33
    12 => "11011111", --  -33
    13 => "11100000", --  -32
    14 => "11100001", --  -31
    15 => "11100011", --  -29
    16 => "11100110", --  -26
    17 => "11101001", --  -23
    18 => "11101101", --  -19
    19 => "11110010", --  -14
    20 => "11111000", --   -8
    21 => "11111110", --   -2
    22 => "00000011", --    3
    23 => "00001001", --    9
    24 => "00001111", --   15
    25 => "00010101", --   21
    26 => "00011010", --   26
    27 => "00011111", --   31
    28 => "00100100", --   36
    29 => "00101000", --   40
    30 => "00101100", --   44
    31 => "00110000", --   48
  );

  constant LUT_1_7_0_DATA : lut_array_t_1 := (
    0 => "00001010", --   10
    1 => "00001011", --   11
    2 => "00001100", --   12
    3 => "00001101", --   13
    4 => "00001110", --   14
    5 => "00001111", --   15
    6 => "00010000", --   16
    7 => "00010000", --   16
    8 => "00010000", --   16
    9 => "00001111", --   15
    10 => "00001111", --   15
    11 => "00001110", --   14
    12 => "00001100", --   12
    13 => "00001010", --   10
    14 => "00001000", --    8
    15 => "00000110", --    6
    16 => "00000100", --    4
    17 => "00000001", --    1
    18 => "11111110", --   -2
    19 => "11111010", --   -6
    20 => "11110111", --   -9
    21 => "11110011", --  -13
    22 => "11101111", --  -17
    23 => "11101011", --  -21
    24 => "11100111", --  -25
    25 => "11100010", --  -30
    26 => "11011110", --  -34
    27 => "11011010", --  -38
    28 => "11010110", --  -42
    29 => "11010010", --  -46
    30 => "11001110", --  -50
    31 => "11001010", --  -54
  );

  constant LUT_1_7_1_DATA : lut_array_t_1 := (
    0 => "00001110", --   14
    1 => "00001110", --   14
    2 => "00001110", --   14
    3 => "00001111", --   15
    4 => "00001111", --   15
    5 => "00010000", --   16
    6 => "00010000", --   16
    7 => "00010000", --   16
    8 => "00010000", --   16
    9 => "00010000", --   16
    10 => "00010000", --   16
    11 => "00001111", --   15
    12 => "00001111", --   15
    13 => "00001101", --   13
    14 => "00001100", --   12
    15 => "00001010", --   10
    16 => "00001000", --    8
    17 => "00000100", --    4
    18 => "00000001", --    1
    19 => "11111101", --   -3
    20 => "11111000", --   -8
    21 => "11110100", --  -12
    22 => "11101110", --  -18
    23 => "11101001", --  -23
    24 => "11100100", --  -28
    25 => "11011110", --  -34
    26 => "11011000", --  -40
    27 => "11010010", --  -46
    28 => "11001100", --  -52
    29 => "11000111", --  -57
    30 => "11000001", --  -63
    31 => "10111100", --  -68
  );

  constant LUT_1_7_2_DATA : lut_array_t_1 := (
    0 => "11100100", --  -28
    1 => "11100101", --  -27
    2 => "11100101", --  -27
    3 => "11100110", --  -26
    4 => "11100111", --  -25
    5 => "11101000", --  -24
    6 => "11101010", --  -22
    7 => "11101011", --  -21
    8 => "11101101", --  -19
    9 => "11101111", --  -17
    10 => "11110001", --  -15
    11 => "11110011", --  -13
    12 => "11110101", --  -11
    13 => "11110111", --   -9
    14 => "11111001", --   -7
    15 => "11111011", --   -5
    16 => "11111110", --   -2
    17 => "00000000", --    0
    18 => "00000011", --    3
    19 => "00000101", --    5
    20 => "00000111", --    7
    21 => "00001010", --   10
    22 => "00001100", --   12
    23 => "00001110", --   14
    24 => "00010000", --   16
    25 => "00010010", --   18
    26 => "00010100", --   20
    27 => "00010101", --   21
    28 => "00010111", --   23
    29 => "00011000", --   24
    30 => "00011001", --   25
    31 => "00011011", --   27
  );

  constant LUT_1_7_3_DATA : lut_array_t_1 := (
    0 => "11111111", --   -1
    1 => "11111111", --   -1
    2 => "11111111", --   -1
    3 => "11111111", --   -1
    4 => "11111111", --   -1
    5 => "00000000", --    0
    6 => "00000000", --    0
    7 => "00000000", --    0
    8 => "00000000", --    0
    9 => "00000000", --    0
    10 => "00000000", --    0
    11 => "00000000", --    0
    12 => "00000000", --    0
    13 => "00000000", --    0
    14 => "00000000", --    0
    15 => "00000000", --    0
    16 => "00000000", --    0
    17 => "00000000", --    0
    18 => "00000001", --    1
    19 => "00000001", --    1
    20 => "00000010", --    2
    21 => "00000011", --    3
    22 => "00000011", --    3
    23 => "00000100", --    4
    24 => "00000101", --    5
    25 => "00000110", --    6
    26 => "00000111", --    7
    27 => "00001000", --    8
    28 => "00001001", --    9
    29 => "00001010", --   10
    30 => "00001011", --   11
    31 => "00001011", --   11
  );

  constant LUT_1_7_4_DATA : lut_array_t_1 := (
    0 => "11100101", --  -27
    1 => "11100100", --  -28
    2 => "11100100", --  -28
    3 => "11100011", --  -29
    4 => "11100100", --  -28
    5 => "11100100", --  -28
    6 => "11100101", --  -27
    7 => "11100110", --  -26
    8 => "11101000", --  -24
    9 => "11101010", --  -22
    10 => "11101100", --  -20
    11 => "11101111", --  -17
    12 => "11110001", --  -15
    13 => "11110100", --  -12
    14 => "11110111", --   -9
    15 => "11111010", --   -6
    16 => "11111101", --   -3
    17 => "11111111", --   -1
    18 => "00000001", --    1
    19 => "00000011", --    3
    20 => "00000101", --    5
    21 => "00000110", --    6
    22 => "00001000", --    8
    23 => "00001001", --    9
    24 => "00001010", --   10
    25 => "00001011", --   11
    26 => "00001100", --   12
    27 => "00001101", --   13
    28 => "00001110", --   14
    29 => "00001111", --   15
    30 => "00001111", --   15
    31 => "00010000", --   16
  );
end package;