library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package PkgLUT is
  -- Layer 0
  subtype lut_output_t_0 is signed(4 downto 0);
  type lut_array_t_0 is array (0 to 63) of lut_output_t_0;


  constant LUT_0_0_0_DATA : lut_array_t_0 := (
    0 => to_signed(2, 5),
    1 => to_signed(3, 5),
    2 => to_signed(3, 5),
    3 => to_signed(3, 5),
    4 => to_signed(3, 5),
    5 => to_signed(3, 5),
    6 => to_signed(3, 5),
    7 => to_signed(3, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(4, 5),
    63 => to_signed(4, 5)
  );

  constant LUT_0_0_1_DATA : lut_array_t_0 := (
    0 => to_signed(3, 5),
    1 => to_signed(3, 5),
    2 => to_signed(3, 5),
    3 => to_signed(3, 5),
    4 => to_signed(3, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(1, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-4, 5),
    15 => to_signed(-4, 5),
    16 => to_signed(-4, 5),
    17 => to_signed(-4, 5),
    18 => to_signed(-4, 5),
    19 => to_signed(-4, 5),
    20 => to_signed(-4, 5),
    21 => to_signed(-4, 5),
    22 => to_signed(-4, 5),
    23 => to_signed(-3, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(2, 5),
    36 => to_signed(3, 5),
    37 => to_signed(3, 5),
    38 => to_signed(3, 5),
    39 => to_signed(4, 5),
    40 => to_signed(4, 5),
    41 => to_signed(4, 5),
    42 => to_signed(5, 5),
    43 => to_signed(5, 5),
    44 => to_signed(5, 5),
    45 => to_signed(6, 5),
    46 => to_signed(6, 5),
    47 => to_signed(6, 5),
    48 => to_signed(7, 5),
    49 => to_signed(7, 5),
    50 => to_signed(8, 5),
    51 => to_signed(8, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(10, 5),
    57 => to_signed(11, 5),
    58 => to_signed(11, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(12, 5),
    62 => to_signed(13, 5),
    63 => to_signed(13, 5)
  );

  constant LUT_0_0_2_DATA : lut_array_t_0 := (
    0 => to_signed(5, 5),
    1 => to_signed(6, 5),
    2 => to_signed(6, 5),
    3 => to_signed(6, 5),
    4 => to_signed(6, 5),
    5 => to_signed(5, 5),
    6 => to_signed(5, 5),
    7 => to_signed(5, 5),
    8 => to_signed(4, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(4, 5),
    20 => to_signed(4, 5),
    21 => to_signed(4, 5),
    22 => to_signed(4, 5),
    23 => to_signed(3, 5),
    24 => to_signed(3, 5),
    25 => to_signed(3, 5),
    26 => to_signed(3, 5),
    27 => to_signed(2, 5),
    28 => to_signed(2, 5),
    29 => to_signed(2, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-3, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-4, 5),
    40 => to_signed(-4, 5),
    41 => to_signed(-5, 5),
    42 => to_signed(-6, 5),
    43 => to_signed(-7, 5),
    44 => to_signed(-7, 5),
    45 => to_signed(-8, 5),
    46 => to_signed(-9, 5),
    47 => to_signed(-10, 5),
    48 => to_signed(-10, 5),
    49 => to_signed(-11, 5),
    50 => to_signed(-12, 5),
    51 => to_signed(-12, 5),
    52 => to_signed(-13, 5),
    53 => to_signed(-14, 5),
    54 => to_signed(-14, 5),
    55 => to_signed(-15, 5),
    56 => to_signed(-15, 5),
    57 => to_signed(-16, 5),
    58 => to_signed(-16, 5),
    59 => to_signed(-16, 5),
    60 => to_signed(-16, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_0_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(2, 5),
    25 => to_signed(2, 5),
    26 => to_signed(2, 5),
    27 => to_signed(2, 5),
    28 => to_signed(2, 5),
    29 => to_signed(2, 5),
    30 => to_signed(2, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-4, 5),
    47 => to_signed(-5, 5),
    48 => to_signed(-5, 5),
    49 => to_signed(-6, 5),
    50 => to_signed(-6, 5),
    51 => to_signed(-7, 5),
    52 => to_signed(-7, 5),
    53 => to_signed(-8, 5),
    54 => to_signed(-8, 5),
    55 => to_signed(-8, 5),
    56 => to_signed(-9, 5),
    57 => to_signed(-9, 5),
    58 => to_signed(-9, 5),
    59 => to_signed(-9, 5),
    60 => to_signed(-9, 5),
    61 => to_signed(-9, 5),
    62 => to_signed(-10, 5),
    63 => to_signed(-10, 5)
  );

  constant LUT_0_0_4_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-3, 5),
    3 => to_signed(-3, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-4, 5),
    6 => to_signed(-4, 5),
    7 => to_signed(-5, 5),
    8 => to_signed(-5, 5),
    9 => to_signed(-6, 5),
    10 => to_signed(-6, 5),
    11 => to_signed(-7, 5),
    12 => to_signed(-7, 5),
    13 => to_signed(-7, 5),
    14 => to_signed(-7, 5),
    15 => to_signed(-8, 5),
    16 => to_signed(-8, 5),
    17 => to_signed(-7, 5),
    18 => to_signed(-7, 5),
    19 => to_signed(-7, 5),
    20 => to_signed(-7, 5),
    21 => to_signed(-6, 5),
    22 => to_signed(-6, 5),
    23 => to_signed(-6, 5),
    24 => to_signed(-5, 5),
    25 => to_signed(-4, 5),
    26 => to_signed(-4, 5),
    27 => to_signed(-3, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(1, 5),
    34 => to_signed(2, 5),
    35 => to_signed(3, 5),
    36 => to_signed(3, 5),
    37 => to_signed(4, 5),
    38 => to_signed(5, 5),
    39 => to_signed(6, 5),
    40 => to_signed(6, 5),
    41 => to_signed(7, 5),
    42 => to_signed(8, 5),
    43 => to_signed(9, 5),
    44 => to_signed(10, 5),
    45 => to_signed(10, 5),
    46 => to_signed(11, 5),
    47 => to_signed(12, 5),
    48 => to_signed(12, 5),
    49 => to_signed(13, 5),
    50 => to_signed(13, 5),
    51 => to_signed(14, 5),
    52 => to_signed(14, 5),
    53 => to_signed(15, 5),
    54 => to_signed(15, 5),
    55 => to_signed(15, 5),
    56 => to_signed(15, 5),
    57 => to_signed(15, 5),
    58 => to_signed(15, 5),
    59 => to_signed(15, 5),
    60 => to_signed(15, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_0_5_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(1, 5),
    60 => to_signed(1, 5),
    61 => to_signed(1, 5),
    62 => to_signed(1, 5),
    63 => to_signed(1, 5)
  );

  constant LUT_0_0_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(0, 5),
    58 => to_signed(0, 5),
    59 => to_signed(0, 5),
    60 => to_signed(0, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_0_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-4, 5),
    53 => to_signed(-4, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-5, 5),
    59 => to_signed(-5, 5),
    60 => to_signed(-5, 5),
    61 => to_signed(-5, 5),
    62 => to_signed(-6, 5),
    63 => to_signed(-6, 5)
  );

  constant LUT_0_1_0_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(4, 5),
    47 => to_signed(5, 5),
    48 => to_signed(5, 5),
    49 => to_signed(5, 5),
    50 => to_signed(6, 5),
    51 => to_signed(6, 5),
    52 => to_signed(6, 5),
    53 => to_signed(6, 5),
    54 => to_signed(7, 5),
    55 => to_signed(7, 5),
    56 => to_signed(7, 5),
    57 => to_signed(8, 5),
    58 => to_signed(8, 5),
    59 => to_signed(8, 5),
    60 => to_signed(8, 5),
    61 => to_signed(9, 5),
    62 => to_signed(9, 5),
    63 => to_signed(10, 5)
  );

  constant LUT_0_1_1_DATA : lut_array_t_0 := (
    0 => to_signed(-5, 5),
    1 => to_signed(-5, 5),
    2 => to_signed(-5, 5),
    3 => to_signed(-5, 5),
    4 => to_signed(-5, 5),
    5 => to_signed(-4, 5),
    6 => to_signed(-4, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-3, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-3, 5),
    21 => to_signed(-3, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(3, 5),
    39 => to_signed(3, 5),
    40 => to_signed(4, 5),
    41 => to_signed(5, 5),
    42 => to_signed(5, 5),
    43 => to_signed(6, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(8, 5),
    47 => to_signed(8, 5),
    48 => to_signed(9, 5),
    49 => to_signed(9, 5),
    50 => to_signed(9, 5),
    51 => to_signed(10, 5),
    52 => to_signed(10, 5),
    53 => to_signed(10, 5),
    54 => to_signed(11, 5),
    55 => to_signed(11, 5),
    56 => to_signed(11, 5),
    57 => to_signed(12, 5),
    58 => to_signed(12, 5),
    59 => to_signed(13, 5),
    60 => to_signed(13, 5),
    61 => to_signed(14, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_1_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-3, 5),
    58 => to_signed(-3, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_1_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(0, 5),
    58 => to_signed(0, 5),
    59 => to_signed(0, 5),
    60 => to_signed(0, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_1_4_DATA : lut_array_t_0 := (
    0 => to_signed(-5, 5),
    1 => to_signed(-5, 5),
    2 => to_signed(-5, 5),
    3 => to_signed(-5, 5),
    4 => to_signed(-5, 5),
    5 => to_signed(-5, 5),
    6 => to_signed(-4, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(2, 5),
    35 => to_signed(2, 5),
    36 => to_signed(3, 5),
    37 => to_signed(3, 5),
    38 => to_signed(3, 5),
    39 => to_signed(3, 5),
    40 => to_signed(4, 5),
    41 => to_signed(4, 5),
    42 => to_signed(4, 5),
    43 => to_signed(4, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(4, 5),
    47 => to_signed(4, 5),
    48 => to_signed(4, 5),
    49 => to_signed(4, 5),
    50 => to_signed(4, 5),
    51 => to_signed(4, 5),
    52 => to_signed(4, 5),
    53 => to_signed(4, 5),
    54 => to_signed(5, 5),
    55 => to_signed(5, 5),
    56 => to_signed(6, 5),
    57 => to_signed(6, 5),
    58 => to_signed(7, 5),
    59 => to_signed(7, 5),
    60 => to_signed(8, 5),
    61 => to_signed(8, 5),
    62 => to_signed(9, 5),
    63 => to_signed(9, 5)
  );

  constant LUT_0_1_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(5, 5),
    47 => to_signed(5, 5),
    48 => to_signed(6, 5),
    49 => to_signed(6, 5),
    50 => to_signed(7, 5),
    51 => to_signed(7, 5),
    52 => to_signed(7, 5),
    53 => to_signed(7, 5),
    54 => to_signed(8, 5),
    55 => to_signed(8, 5),
    56 => to_signed(8, 5),
    57 => to_signed(8, 5),
    58 => to_signed(8, 5),
    59 => to_signed(8, 5),
    60 => to_signed(8, 5),
    61 => to_signed(9, 5),
    62 => to_signed(9, 5),
    63 => to_signed(9, 5)
  );

  constant LUT_0_1_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(0, 5),
    58 => to_signed(0, 5),
    59 => to_signed(0, 5),
    60 => to_signed(0, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_1_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(4, 5),
    53 => to_signed(4, 5),
    54 => to_signed(4, 5),
    55 => to_signed(4, 5),
    56 => to_signed(5, 5),
    57 => to_signed(5, 5),
    58 => to_signed(5, 5),
    59 => to_signed(5, 5),
    60 => to_signed(5, 5),
    61 => to_signed(6, 5),
    62 => to_signed(6, 5),
    63 => to_signed(6, 5)
  );

  constant LUT_0_2_0_DATA : lut_array_t_0 := (
    0 => to_signed(2, 5),
    1 => to_signed(2, 5),
    2 => to_signed(3, 5),
    3 => to_signed(3, 5),
    4 => to_signed(3, 5),
    5 => to_signed(3, 5),
    6 => to_signed(4, 5),
    7 => to_signed(4, 5),
    8 => to_signed(4, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(5, 5),
    12 => to_signed(5, 5),
    13 => to_signed(5, 5),
    14 => to_signed(4, 5),
    15 => to_signed(4, 5),
    16 => to_signed(4, 5),
    17 => to_signed(4, 5),
    18 => to_signed(3, 5),
    19 => to_signed(3, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(0, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-2, 5),
    32 => to_signed(-2, 5),
    33 => to_signed(-2, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-3, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-4, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-4, 5),
    47 => to_signed(-4, 5),
    48 => to_signed(-5, 5),
    49 => to_signed(-5, 5),
    50 => to_signed(-5, 5),
    51 => to_signed(-6, 5),
    52 => to_signed(-6, 5),
    53 => to_signed(-7, 5),
    54 => to_signed(-7, 5),
    55 => to_signed(-8, 5),
    56 => to_signed(-8, 5),
    57 => to_signed(-9, 5),
    58 => to_signed(-9, 5),
    59 => to_signed(-10, 5),
    60 => to_signed(-10, 5),
    61 => to_signed(-10, 5),
    62 => to_signed(-10, 5),
    63 => to_signed(-10, 5)
  );

  constant LUT_0_2_1_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(3, 5),
    9 => to_signed(3, 5),
    10 => to_signed(3, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(3, 5),
    20 => to_signed(3, 5),
    21 => to_signed(3, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(2, 5),
    25 => to_signed(2, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-4, 5),
    44 => to_signed(-5, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-6, 5),
    47 => to_signed(-7, 5),
    48 => to_signed(-7, 5),
    49 => to_signed(-8, 5),
    50 => to_signed(-9, 5),
    51 => to_signed(-9, 5),
    52 => to_signed(-10, 5),
    53 => to_signed(-11, 5),
    54 => to_signed(-12, 5),
    55 => to_signed(-12, 5),
    56 => to_signed(-13, 5),
    57 => to_signed(-14, 5),
    58 => to_signed(-14, 5),
    59 => to_signed(-15, 5),
    60 => to_signed(-15, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_2_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(2, 5),
    25 => to_signed(2, 5),
    26 => to_signed(2, 5),
    27 => to_signed(2, 5),
    28 => to_signed(2, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-4, 5),
    41 => to_signed(-4, 5),
    42 => to_signed(-5, 5),
    43 => to_signed(-5, 5),
    44 => to_signed(-5, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-5, 5),
    47 => to_signed(-6, 5),
    48 => to_signed(-6, 5),
    49 => to_signed(-6, 5),
    50 => to_signed(-6, 5),
    51 => to_signed(-6, 5),
    52 => to_signed(-6, 5),
    53 => to_signed(-6, 5),
    54 => to_signed(-6, 5),
    55 => to_signed(-7, 5),
    56 => to_signed(-7, 5),
    57 => to_signed(-7, 5),
    58 => to_signed(-8, 5),
    59 => to_signed(-8, 5),
    60 => to_signed(-9, 5),
    61 => to_signed(-9, 5),
    62 => to_signed(-9, 5),
    63 => to_signed(-10, 5)
  );

  constant LUT_0_2_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(3, 5),
    46 => to_signed(3, 5),
    47 => to_signed(4, 5),
    48 => to_signed(4, 5),
    49 => to_signed(4, 5),
    50 => to_signed(5, 5),
    51 => to_signed(5, 5),
    52 => to_signed(5, 5),
    53 => to_signed(6, 5),
    54 => to_signed(6, 5),
    55 => to_signed(6, 5),
    56 => to_signed(6, 5),
    57 => to_signed(7, 5),
    58 => to_signed(7, 5),
    59 => to_signed(7, 5),
    60 => to_signed(7, 5),
    61 => to_signed(7, 5),
    62 => to_signed(7, 5),
    63 => to_signed(7, 5)
  );

  constant LUT_0_2_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(2, 5),
    63 => to_signed(2, 5)
  );

  constant LUT_0_2_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(3, 5),
    41 => to_signed(3, 5),
    42 => to_signed(4, 5),
    43 => to_signed(4, 5),
    44 => to_signed(5, 5),
    45 => to_signed(5, 5),
    46 => to_signed(6, 5),
    47 => to_signed(6, 5),
    48 => to_signed(6, 5),
    49 => to_signed(7, 5),
    50 => to_signed(7, 5),
    51 => to_signed(8, 5),
    52 => to_signed(8, 5),
    53 => to_signed(8, 5),
    54 => to_signed(9, 5),
    55 => to_signed(9, 5),
    56 => to_signed(10, 5),
    57 => to_signed(11, 5),
    58 => to_signed(11, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(13, 5),
    62 => to_signed(14, 5),
    63 => to_signed(14, 5)
  );

  constant LUT_0_2_6_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-5, 5),
    10 => to_signed(-6, 5),
    11 => to_signed(-6, 5),
    12 => to_signed(-6, 5),
    13 => to_signed(-7, 5),
    14 => to_signed(-7, 5),
    15 => to_signed(-6, 5),
    16 => to_signed(-6, 5),
    17 => to_signed(-6, 5),
    18 => to_signed(-6, 5),
    19 => to_signed(-5, 5),
    20 => to_signed(-5, 5),
    21 => to_signed(-4, 5),
    22 => to_signed(-4, 5),
    23 => to_signed(-4, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(3, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(5, 5),
    47 => to_signed(5, 5),
    48 => to_signed(6, 5),
    49 => to_signed(6, 5),
    50 => to_signed(7, 5),
    51 => to_signed(8, 5),
    52 => to_signed(8, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(11, 5),
    57 => to_signed(11, 5),
    58 => to_signed(11, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(12, 5),
    62 => to_signed(12, 5),
    63 => to_signed(12, 5)
  );

  constant LUT_0_2_7_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-3, 5),
    3 => to_signed(-3, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-4, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-4, 5),
    12 => to_signed(-4, 5),
    13 => to_signed(-4, 5),
    14 => to_signed(-4, 5),
    15 => to_signed(-4, 5),
    16 => to_signed(-4, 5),
    17 => to_signed(-4, 5),
    18 => to_signed(-4, 5),
    19 => to_signed(-4, 5),
    20 => to_signed(-4, 5),
    21 => to_signed(-3, 5),
    22 => to_signed(-3, 5),
    23 => to_signed(-3, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(2, 5),
    36 => to_signed(2, 5),
    37 => to_signed(3, 5),
    38 => to_signed(3, 5),
    39 => to_signed(4, 5),
    40 => to_signed(4, 5),
    41 => to_signed(5, 5),
    42 => to_signed(5, 5),
    43 => to_signed(6, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(8, 5),
    47 => to_signed(9, 5),
    48 => to_signed(9, 5),
    49 => to_signed(10, 5),
    50 => to_signed(11, 5),
    51 => to_signed(11, 5),
    52 => to_signed(12, 5),
    53 => to_signed(12, 5),
    54 => to_signed(13, 5),
    55 => to_signed(13, 5),
    56 => to_signed(14, 5),
    57 => to_signed(14, 5),
    58 => to_signed(15, 5),
    59 => to_signed(15, 5),
    60 => to_signed(15, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_3_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-3, 5),
    27 => to_signed(-3, 5),
    28 => to_signed(-3, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(3, 5),
    47 => to_signed(3, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_3_1_DATA : lut_array_t_0 := (
    0 => to_signed(2, 5),
    1 => to_signed(3, 5),
    2 => to_signed(3, 5),
    3 => to_signed(3, 5),
    4 => to_signed(4, 5),
    5 => to_signed(4, 5),
    6 => to_signed(4, 5),
    7 => to_signed(5, 5),
    8 => to_signed(5, 5),
    9 => to_signed(5, 5),
    10 => to_signed(6, 5),
    11 => to_signed(6, 5),
    12 => to_signed(6, 5),
    13 => to_signed(6, 5),
    14 => to_signed(6, 5),
    15 => to_signed(7, 5),
    16 => to_signed(7, 5),
    17 => to_signed(7, 5),
    18 => to_signed(7, 5),
    19 => to_signed(7, 5),
    20 => to_signed(7, 5),
    21 => to_signed(7, 5),
    22 => to_signed(7, 5),
    23 => to_signed(6, 5),
    24 => to_signed(6, 5),
    25 => to_signed(5, 5),
    26 => to_signed(5, 5),
    27 => to_signed(4, 5),
    28 => to_signed(2, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-2, 5),
    33 => to_signed(-4, 5),
    34 => to_signed(-5, 5),
    35 => to_signed(-6, 5),
    36 => to_signed(-7, 5),
    37 => to_signed(-7, 5),
    38 => to_signed(-8, 5),
    39 => to_signed(-9, 5),
    40 => to_signed(-9, 5),
    41 => to_signed(-9, 5),
    42 => to_signed(-9, 5),
    43 => to_signed(-9, 5),
    44 => to_signed(-9, 5),
    45 => to_signed(-9, 5),
    46 => to_signed(-9, 5),
    47 => to_signed(-9, 5),
    48 => to_signed(-9, 5),
    49 => to_signed(-9, 5),
    50 => to_signed(-9, 5),
    51 => to_signed(-10, 5),
    52 => to_signed(-10, 5),
    53 => to_signed(-10, 5),
    54 => to_signed(-11, 5),
    55 => to_signed(-11, 5),
    56 => to_signed(-12, 5),
    57 => to_signed(-13, 5),
    58 => to_signed(-13, 5),
    59 => to_signed(-14, 5),
    60 => to_signed(-15, 5),
    61 => to_signed(-15, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_3_2_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-3, 5),
    57 => to_signed(-3, 5),
    58 => to_signed(-3, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_3_3_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(2, 5),
    37 => to_signed(3, 5),
    38 => to_signed(3, 5),
    39 => to_signed(4, 5),
    40 => to_signed(5, 5),
    41 => to_signed(5, 5),
    42 => to_signed(6, 5),
    43 => to_signed(7, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(8, 5),
    47 => to_signed(8, 5),
    48 => to_signed(8, 5),
    49 => to_signed(8, 5),
    50 => to_signed(8, 5),
    51 => to_signed(9, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(11, 5),
    57 => to_signed(11, 5),
    58 => to_signed(12, 5),
    59 => to_signed(12, 5),
    60 => to_signed(13, 5),
    61 => to_signed(14, 5),
    62 => to_signed(14, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_3_4_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(3, 5),
    41 => to_signed(4, 5),
    42 => to_signed(5, 5),
    43 => to_signed(6, 5),
    44 => to_signed(7, 5),
    45 => to_signed(8, 5),
    46 => to_signed(9, 5),
    47 => to_signed(9, 5),
    48 => to_signed(10, 5),
    49 => to_signed(10, 5),
    50 => to_signed(10, 5),
    51 => to_signed(11, 5),
    52 => to_signed(11, 5),
    53 => to_signed(11, 5),
    54 => to_signed(12, 5),
    55 => to_signed(12, 5),
    56 => to_signed(12, 5),
    57 => to_signed(13, 5),
    58 => to_signed(13, 5),
    59 => to_signed(13, 5),
    60 => to_signed(14, 5),
    61 => to_signed(14, 5),
    62 => to_signed(14, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_3_5_DATA : lut_array_t_0 := (
    0 => to_signed(4, 5),
    1 => to_signed(5, 5),
    2 => to_signed(5, 5),
    3 => to_signed(6, 5),
    4 => to_signed(7, 5),
    5 => to_signed(8, 5),
    6 => to_signed(9, 5),
    7 => to_signed(9, 5),
    8 => to_signed(10, 5),
    9 => to_signed(10, 5),
    10 => to_signed(11, 5),
    11 => to_signed(11, 5),
    12 => to_signed(11, 5),
    13 => to_signed(11, 5),
    14 => to_signed(11, 5),
    15 => to_signed(11, 5),
    16 => to_signed(11, 5),
    17 => to_signed(10, 5),
    18 => to_signed(10, 5),
    19 => to_signed(10, 5),
    20 => to_signed(9, 5),
    21 => to_signed(9, 5),
    22 => to_signed(8, 5),
    23 => to_signed(7, 5),
    24 => to_signed(7, 5),
    25 => to_signed(6, 5),
    26 => to_signed(4, 5),
    27 => to_signed(3, 5),
    28 => to_signed(2, 5),
    29 => to_signed(0, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-3, 5),
    32 => to_signed(-4, 5),
    33 => to_signed(-6, 5),
    34 => to_signed(-7, 5),
    35 => to_signed(-8, 5),
    36 => to_signed(-9, 5),
    37 => to_signed(-9, 5),
    38 => to_signed(-10, 5),
    39 => to_signed(-11, 5),
    40 => to_signed(-12, 5),
    41 => to_signed(-13, 5),
    42 => to_signed(-14, 5),
    43 => to_signed(-14, 5),
    44 => to_signed(-15, 5),
    45 => to_signed(-16, 5),
    46 => to_signed(-16, 5),
    47 => to_signed(-16, 5),
    48 => to_signed(-16, 5),
    49 => to_signed(-16, 5),
    50 => to_signed(-16, 5),
    51 => to_signed(-16, 5),
    52 => to_signed(-16, 5),
    53 => to_signed(-16, 5),
    54 => to_signed(-16, 5),
    55 => to_signed(-16, 5),
    56 => to_signed(-16, 5),
    57 => to_signed(-16, 5),
    58 => to_signed(-16, 5),
    59 => to_signed(-16, 5),
    60 => to_signed(-16, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_3_6_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-3, 5),
    2 => to_signed(-3, 5),
    3 => to_signed(-4, 5),
    4 => to_signed(-5, 5),
    5 => to_signed(-6, 5),
    6 => to_signed(-7, 5),
    7 => to_signed(-8, 5),
    8 => to_signed(-9, 5),
    9 => to_signed(-11, 5),
    10 => to_signed(-12, 5),
    11 => to_signed(-13, 5),
    12 => to_signed(-14, 5),
    13 => to_signed(-15, 5),
    14 => to_signed(-16, 5),
    15 => to_signed(-16, 5),
    16 => to_signed(-16, 5),
    17 => to_signed(-16, 5),
    18 => to_signed(-16, 5),
    19 => to_signed(-16, 5),
    20 => to_signed(-16, 5),
    21 => to_signed(-15, 5),
    22 => to_signed(-14, 5),
    23 => to_signed(-13, 5),
    24 => to_signed(-12, 5),
    25 => to_signed(-10, 5),
    26 => to_signed(-8, 5),
    27 => to_signed(-6, 5),
    28 => to_signed(-4, 5),
    29 => to_signed(-3, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(3, 5),
    33 => to_signed(4, 5),
    34 => to_signed(5, 5),
    35 => to_signed(7, 5),
    36 => to_signed(8, 5),
    37 => to_signed(9, 5),
    38 => to_signed(9, 5),
    39 => to_signed(10, 5),
    40 => to_signed(11, 5),
    41 => to_signed(12, 5),
    42 => to_signed(12, 5),
    43 => to_signed(13, 5),
    44 => to_signed(14, 5),
    45 => to_signed(14, 5),
    46 => to_signed(15, 5),
    47 => to_signed(15, 5),
    48 => to_signed(15, 5),
    49 => to_signed(15, 5),
    50 => to_signed(15, 5),
    51 => to_signed(15, 5),
    52 => to_signed(15, 5),
    53 => to_signed(15, 5),
    54 => to_signed(15, 5),
    55 => to_signed(15, 5),
    56 => to_signed(15, 5),
    57 => to_signed(15, 5),
    58 => to_signed(15, 5),
    59 => to_signed(15, 5),
    60 => to_signed(15, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_3_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-3, 5),
    10 => to_signed(-3, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-4, 5),
    15 => to_signed(-4, 5),
    16 => to_signed(-4, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-3, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(0, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(2, 5),
    26 => to_signed(3, 5),
    27 => to_signed(3, 5),
    28 => to_signed(3, 5),
    29 => to_signed(3, 5),
    30 => to_signed(3, 5),
    31 => to_signed(3, 5),
    32 => to_signed(3, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(0, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-4, 5),
    50 => to_signed(-4, 5),
    51 => to_signed(-4, 5),
    52 => to_signed(-4, 5),
    53 => to_signed(-4, 5),
    54 => to_signed(-5, 5),
    55 => to_signed(-5, 5),
    56 => to_signed(-5, 5),
    57 => to_signed(-6, 5),
    58 => to_signed(-6, 5),
    59 => to_signed(-7, 5),
    60 => to_signed(-7, 5),
    61 => to_signed(-8, 5),
    62 => to_signed(-8, 5),
    63 => to_signed(-9, 5)
  );

  constant LUT_0_4_0_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(3, 5),
    8 => to_signed(3, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(5, 5),
    12 => to_signed(5, 5),
    13 => to_signed(6, 5),
    14 => to_signed(6, 5),
    15 => to_signed(6, 5),
    16 => to_signed(6, 5),
    17 => to_signed(5, 5),
    18 => to_signed(5, 5),
    19 => to_signed(4, 5),
    20 => to_signed(3, 5),
    21 => to_signed(3, 5),
    22 => to_signed(2, 5),
    23 => to_signed(1, 5),
    24 => to_signed(0, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-3, 5),
    30 => to_signed(-3, 5),
    31 => to_signed(-3, 5),
    32 => to_signed(-3, 5),
    33 => to_signed(-3, 5),
    34 => to_signed(-3, 5),
    35 => to_signed(-3, 5),
    36 => to_signed(-3, 5),
    37 => to_signed(-3, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-4, 5),
    44 => to_signed(-4, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-4, 5),
    47 => to_signed(-4, 5),
    48 => to_signed(-4, 5),
    49 => to_signed(-4, 5),
    50 => to_signed(-5, 5),
    51 => to_signed(-5, 5),
    52 => to_signed(-5, 5),
    53 => to_signed(-5, 5),
    54 => to_signed(-6, 5),
    55 => to_signed(-6, 5),
    56 => to_signed(-6, 5),
    57 => to_signed(-6, 5),
    58 => to_signed(-7, 5),
    59 => to_signed(-7, 5),
    60 => to_signed(-7, 5),
    61 => to_signed(-7, 5),
    62 => to_signed(-7, 5),
    63 => to_signed(-7, 5)
  );

  constant LUT_0_4_1_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(3, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(5, 5),
    47 => to_signed(5, 5),
    48 => to_signed(5, 5),
    49 => to_signed(6, 5),
    50 => to_signed(6, 5),
    51 => to_signed(6, 5),
    52 => to_signed(6, 5),
    53 => to_signed(6, 5),
    54 => to_signed(6, 5),
    55 => to_signed(6, 5),
    56 => to_signed(6, 5),
    57 => to_signed(6, 5),
    58 => to_signed(6, 5),
    59 => to_signed(6, 5),
    60 => to_signed(6, 5),
    61 => to_signed(6, 5),
    62 => to_signed(6, 5),
    63 => to_signed(6, 5)
  );

  constant LUT_0_4_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(3, 5),
    20 => to_signed(3, 5),
    21 => to_signed(3, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(2, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-4, 5),
    41 => to_signed(-4, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-5, 5),
    44 => to_signed(-5, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-5, 5),
    47 => to_signed(-6, 5),
    48 => to_signed(-6, 5),
    49 => to_signed(-6, 5),
    50 => to_signed(-6, 5),
    51 => to_signed(-7, 5),
    52 => to_signed(-7, 5),
    53 => to_signed(-7, 5),
    54 => to_signed(-8, 5),
    55 => to_signed(-8, 5),
    56 => to_signed(-8, 5),
    57 => to_signed(-9, 5),
    58 => to_signed(-9, 5),
    59 => to_signed(-10, 5),
    60 => to_signed(-10, 5),
    61 => to_signed(-11, 5),
    62 => to_signed(-11, 5),
    63 => to_signed(-12, 5)
  );

  constant LUT_0_4_3_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(3, 5),
    10 => to_signed(3, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(3, 5),
    20 => to_signed(3, 5),
    21 => to_signed(3, 5),
    22 => to_signed(3, 5),
    23 => to_signed(2, 5),
    24 => to_signed(2, 5),
    25 => to_signed(2, 5),
    26 => to_signed(2, 5),
    27 => to_signed(2, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-4, 5),
    41 => to_signed(-5, 5),
    42 => to_signed(-5, 5),
    43 => to_signed(-6, 5),
    44 => to_signed(-7, 5),
    45 => to_signed(-7, 5),
    46 => to_signed(-8, 5),
    47 => to_signed(-9, 5),
    48 => to_signed(-9, 5),
    49 => to_signed(-10, 5),
    50 => to_signed(-10, 5),
    51 => to_signed(-10, 5),
    52 => to_signed(-10, 5),
    53 => to_signed(-11, 5),
    54 => to_signed(-11, 5),
    55 => to_signed(-11, 5),
    56 => to_signed(-11, 5),
    57 => to_signed(-11, 5),
    58 => to_signed(-11, 5),
    59 => to_signed(-11, 5),
    60 => to_signed(-11, 5),
    61 => to_signed(-12, 5),
    62 => to_signed(-12, 5),
    63 => to_signed(-12, 5)
  );

  constant LUT_0_4_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_4_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(3, 5),
    42 => to_signed(3, 5),
    43 => to_signed(4, 5),
    44 => to_signed(4, 5),
    45 => to_signed(5, 5),
    46 => to_signed(5, 5),
    47 => to_signed(6, 5),
    48 => to_signed(6, 5),
    49 => to_signed(6, 5),
    50 => to_signed(7, 5),
    51 => to_signed(7, 5),
    52 => to_signed(7, 5),
    53 => to_signed(7, 5),
    54 => to_signed(8, 5),
    55 => to_signed(8, 5),
    56 => to_signed(8, 5),
    57 => to_signed(9, 5),
    58 => to_signed(9, 5),
    59 => to_signed(9, 5),
    60 => to_signed(10, 5),
    61 => to_signed(10, 5),
    62 => to_signed(11, 5),
    63 => to_signed(11, 5)
  );

  constant LUT_0_4_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-3, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-4, 5),
    14 => to_signed(-4, 5),
    15 => to_signed(-4, 5),
    16 => to_signed(-4, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-3, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-3, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(2, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(4, 5),
    60 => to_signed(5, 5),
    61 => to_signed(5, 5),
    62 => to_signed(5, 5),
    63 => to_signed(6, 5)
  );

  constant LUT_0_4_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-2, 5),
    14 => to_signed(-2, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(3, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(4, 5),
    51 => to_signed(4, 5),
    52 => to_signed(5, 5),
    53 => to_signed(5, 5),
    54 => to_signed(5, 5),
    55 => to_signed(6, 5),
    56 => to_signed(6, 5),
    57 => to_signed(7, 5),
    58 => to_signed(7, 5),
    59 => to_signed(8, 5),
    60 => to_signed(8, 5),
    61 => to_signed(8, 5),
    62 => to_signed(8, 5),
    63 => to_signed(8, 5)
  );

  constant LUT_0_5_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(0, 5),
    54 => to_signed(0, 5),
    55 => to_signed(0, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(0, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_5_1_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(4, 5),
    45 => to_signed(4, 5),
    46 => to_signed(4, 5),
    47 => to_signed(5, 5),
    48 => to_signed(5, 5),
    49 => to_signed(5, 5),
    50 => to_signed(5, 5),
    51 => to_signed(5, 5),
    52 => to_signed(6, 5),
    53 => to_signed(6, 5),
    54 => to_signed(6, 5),
    55 => to_signed(6, 5),
    56 => to_signed(6, 5),
    57 => to_signed(6, 5),
    58 => to_signed(7, 5),
    59 => to_signed(7, 5),
    60 => to_signed(7, 5),
    61 => to_signed(7, 5),
    62 => to_signed(7, 5),
    63 => to_signed(8, 5)
  );

  constant LUT_0_5_2_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_5_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(1, 5),
    57 => to_signed(1, 5),
    58 => to_signed(1, 5),
    59 => to_signed(1, 5),
    60 => to_signed(1, 5),
    61 => to_signed(1, 5),
    62 => to_signed(1, 5),
    63 => to_signed(1, 5)
  );

  constant LUT_0_5_4_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-3, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-3, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(2, 5),
    32 => to_signed(2, 5),
    33 => to_signed(2, 5),
    34 => to_signed(3, 5),
    35 => to_signed(3, 5),
    36 => to_signed(3, 5),
    37 => to_signed(4, 5),
    38 => to_signed(4, 5),
    39 => to_signed(5, 5),
    40 => to_signed(5, 5),
    41 => to_signed(6, 5),
    42 => to_signed(6, 5),
    43 => to_signed(7, 5),
    44 => to_signed(7, 5),
    45 => to_signed(8, 5),
    46 => to_signed(8, 5),
    47 => to_signed(9, 5),
    48 => to_signed(10, 5),
    49 => to_signed(10, 5),
    50 => to_signed(11, 5),
    51 => to_signed(11, 5),
    52 => to_signed(12, 5),
    53 => to_signed(12, 5),
    54 => to_signed(13, 5),
    55 => to_signed(13, 5),
    56 => to_signed(14, 5),
    57 => to_signed(15, 5),
    58 => to_signed(15, 5),
    59 => to_signed(15, 5),
    60 => to_signed(15, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_5_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-4, 5),
    6 => to_signed(-6, 5),
    7 => to_signed(-7, 5),
    8 => to_signed(-9, 5),
    9 => to_signed(-10, 5),
    10 => to_signed(-11, 5),
    11 => to_signed(-12, 5),
    12 => to_signed(-13, 5),
    13 => to_signed(-12, 5),
    14 => to_signed(-12, 5),
    15 => to_signed(-10, 5),
    16 => to_signed(-9, 5),
    17 => to_signed(-7, 5),
    18 => to_signed(-5, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(0, 5),
    22 => to_signed(1, 5),
    23 => to_signed(2, 5),
    24 => to_signed(3, 5),
    25 => to_signed(3, 5),
    26 => to_signed(4, 5),
    27 => to_signed(4, 5),
    28 => to_signed(4, 5),
    29 => to_signed(3, 5),
    30 => to_signed(3, 5),
    31 => to_signed(3, 5),
    32 => to_signed(2, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(2, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_5_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(3, 5),
    45 => to_signed(3, 5),
    46 => to_signed(3, 5),
    47 => to_signed(4, 5),
    48 => to_signed(4, 5),
    49 => to_signed(4, 5),
    50 => to_signed(4, 5),
    51 => to_signed(4, 5),
    52 => to_signed(5, 5),
    53 => to_signed(5, 5),
    54 => to_signed(5, 5),
    55 => to_signed(5, 5),
    56 => to_signed(5, 5),
    57 => to_signed(6, 5),
    58 => to_signed(6, 5),
    59 => to_signed(6, 5),
    60 => to_signed(6, 5),
    61 => to_signed(7, 5),
    62 => to_signed(7, 5),
    63 => to_signed(7, 5)
  );

  constant LUT_0_5_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(3, 5),
    45 => to_signed(4, 5),
    46 => to_signed(4, 5),
    47 => to_signed(4, 5),
    48 => to_signed(5, 5),
    49 => to_signed(5, 5),
    50 => to_signed(5, 5),
    51 => to_signed(6, 5),
    52 => to_signed(6, 5),
    53 => to_signed(7, 5),
    54 => to_signed(7, 5),
    55 => to_signed(7, 5),
    56 => to_signed(8, 5),
    57 => to_signed(8, 5),
    58 => to_signed(8, 5),
    59 => to_signed(9, 5),
    60 => to_signed(9, 5),
    61 => to_signed(9, 5),
    62 => to_signed(9, 5),
    63 => to_signed(9, 5)
  );

  constant LUT_0_6_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(0, 5),
    54 => to_signed(0, 5),
    55 => to_signed(0, 5),
    56 => to_signed(0, 5),
    57 => to_signed(0, 5),
    58 => to_signed(0, 5),
    59 => to_signed(0, 5),
    60 => to_signed(0, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_6_1_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_6_2_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_6_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_6_4_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-4, 5),
    53 => to_signed(-4, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-5, 5),
    58 => to_signed(-5, 5),
    59 => to_signed(-5, 5),
    60 => to_signed(-6, 5),
    61 => to_signed(-6, 5),
    62 => to_signed(-6, 5),
    63 => to_signed(-7, 5)
  );

  constant LUT_0_6_5_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_6_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(0, 5),
    54 => to_signed(0, 5),
    55 => to_signed(1, 5),
    56 => to_signed(1, 5),
    57 => to_signed(1, 5),
    58 => to_signed(1, 5),
    59 => to_signed(1, 5),
    60 => to_signed(1, 5),
    61 => to_signed(1, 5),
    62 => to_signed(1, 5),
    63 => to_signed(1, 5)
  );

  constant LUT_0_6_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_7_0_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-3, 5),
    8 => to_signed(-3, 5),
    9 => to_signed(-3, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-4, 5),
    12 => to_signed(-4, 5),
    13 => to_signed(-4, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(3, 5),
    47 => to_signed(3, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(4, 5),
    54 => to_signed(4, 5),
    55 => to_signed(4, 5),
    56 => to_signed(4, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(4, 5),
    60 => to_signed(5, 5),
    61 => to_signed(5, 5),
    62 => to_signed(5, 5),
    63 => to_signed(5, 5)
  );

  constant LUT_0_7_1_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_7_2_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-2, 5),
    14 => to_signed(-2, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_7_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-2, 5),
    14 => to_signed(-2, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(3, 5),
    45 => to_signed(3, 5),
    46 => to_signed(3, 5),
    47 => to_signed(3, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(4, 5),
    55 => to_signed(4, 5),
    56 => to_signed(4, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(4, 5),
    60 => to_signed(4, 5),
    61 => to_signed(4, 5),
    62 => to_signed(5, 5),
    63 => to_signed(5, 5)
  );

  constant LUT_0_7_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-2, 5),
    14 => to_signed(-2, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(4, 5),
    62 => to_signed(4, 5),
    63 => to_signed(4, 5)
  );

  constant LUT_0_7_5_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(2, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(3, 5),
    5 => to_signed(3, 5),
    6 => to_signed(3, 5),
    7 => to_signed(3, 5),
    8 => to_signed(4, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-3, 5),
    32 => to_signed(-3, 5),
    33 => to_signed(-3, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_7_6_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-3, 5),
    10 => to_signed(-3, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-2, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(2, 5),
    29 => to_signed(2, 5),
    30 => to_signed(2, 5),
    31 => to_signed(2, 5),
    32 => to_signed(2, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(2, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(3, 5),
    49 => to_signed(3, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_7_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(2, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_8_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_8_1_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_8_2_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_8_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-4, 5),
    59 => to_signed(-5, 5),
    60 => to_signed(-5, 5),
    61 => to_signed(-5, 5),
    62 => to_signed(-5, 5),
    63 => to_signed(-5, 5)
  );

  constant LUT_0_8_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_8_5_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(2, 5),
    63 => to_signed(2, 5)
  );

  constant LUT_0_8_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_8_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-1, 5)
  );

  constant LUT_0_9_0_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(4, 5),
    63 => to_signed(4, 5)
  );

  constant LUT_0_9_1_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_9_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_9_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-4, 5),
    53 => to_signed(-4, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-5, 5),
    58 => to_signed(-5, 5),
    59 => to_signed(-5, 5),
    60 => to_signed(-5, 5),
    61 => to_signed(-6, 5),
    62 => to_signed(-6, 5),
    63 => to_signed(-6, 5)
  );

  constant LUT_0_9_4_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(2, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(3, 5),
    44 => to_signed(3, 5),
    45 => to_signed(3, 5),
    46 => to_signed(4, 5),
    47 => to_signed(4, 5),
    48 => to_signed(4, 5),
    49 => to_signed(5, 5),
    50 => to_signed(5, 5),
    51 => to_signed(5, 5),
    52 => to_signed(6, 5),
    53 => to_signed(6, 5),
    54 => to_signed(6, 5),
    55 => to_signed(7, 5),
    56 => to_signed(7, 5),
    57 => to_signed(7, 5),
    58 => to_signed(8, 5),
    59 => to_signed(8, 5),
    60 => to_signed(9, 5),
    61 => to_signed(9, 5),
    62 => to_signed(9, 5),
    63 => to_signed(10, 5)
  );

  constant LUT_0_9_5_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-4, 5),
    59 => to_signed(-4, 5),
    60 => to_signed(-4, 5),
    61 => to_signed(-5, 5),
    62 => to_signed(-5, 5),
    63 => to_signed(-5, 5)
  );

  constant LUT_0_9_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_9_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(2, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(4, 5),
    60 => to_signed(4, 5),
    61 => to_signed(4, 5),
    62 => to_signed(5, 5),
    63 => to_signed(5, 5)
  );

  constant LUT_0_10_0_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_10_1_DATA : lut_array_t_0 := (
    0 => to_signed(-5, 5),
    1 => to_signed(-5, 5),
    2 => to_signed(-5, 5),
    3 => to_signed(-6, 5),
    4 => to_signed(-6, 5),
    5 => to_signed(-6, 5),
    6 => to_signed(-6, 5),
    7 => to_signed(-6, 5),
    8 => to_signed(-6, 5),
    9 => to_signed(-6, 5),
    10 => to_signed(-5, 5),
    11 => to_signed(-5, 5),
    12 => to_signed(-5, 5),
    13 => to_signed(-4, 5),
    14 => to_signed(-4, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(2, 5),
    36 => to_signed(3, 5),
    37 => to_signed(3, 5),
    38 => to_signed(3, 5),
    39 => to_signed(4, 5),
    40 => to_signed(4, 5),
    41 => to_signed(4, 5),
    42 => to_signed(4, 5),
    43 => to_signed(5, 5),
    44 => to_signed(5, 5),
    45 => to_signed(5, 5),
    46 => to_signed(5, 5),
    47 => to_signed(6, 5),
    48 => to_signed(6, 5),
    49 => to_signed(6, 5),
    50 => to_signed(7, 5),
    51 => to_signed(7, 5),
    52 => to_signed(7, 5),
    53 => to_signed(8, 5),
    54 => to_signed(8, 5),
    55 => to_signed(9, 5),
    56 => to_signed(9, 5),
    57 => to_signed(9, 5),
    58 => to_signed(10, 5),
    59 => to_signed(10, 5),
    60 => to_signed(11, 5),
    61 => to_signed(11, 5),
    62 => to_signed(11, 5),
    63 => to_signed(12, 5)
  );

  constant LUT_0_10_2_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(2, 5),
    63 => to_signed(2, 5)
  );

  constant LUT_0_10_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-3, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-4, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-4, 5),
    47 => to_signed(-4, 5),
    48 => to_signed(-5, 5),
    49 => to_signed(-5, 5),
    50 => to_signed(-5, 5),
    51 => to_signed(-5, 5),
    52 => to_signed(-6, 5),
    53 => to_signed(-6, 5),
    54 => to_signed(-6, 5),
    55 => to_signed(-7, 5),
    56 => to_signed(-7, 5),
    57 => to_signed(-7, 5),
    58 => to_signed(-8, 5),
    59 => to_signed(-8, 5),
    60 => to_signed(-8, 5),
    61 => to_signed(-9, 5),
    62 => to_signed(-9, 5),
    63 => to_signed(-10, 5)
  );

  constant LUT_0_10_4_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(2, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(3, 5),
    51 => to_signed(3, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(4, 5),
    56 => to_signed(4, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(5, 5),
    60 => to_signed(5, 5),
    61 => to_signed(5, 5),
    62 => to_signed(5, 5),
    63 => to_signed(5, 5)
  );

  constant LUT_0_10_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(4, 5),
    62 => to_signed(4, 5),
    63 => to_signed(4, 5)
  );

  constant LUT_0_10_6_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(2, 5),
    2 => to_signed(2, 5),
    3 => to_signed(3, 5),
    4 => to_signed(3, 5),
    5 => to_signed(4, 5),
    6 => to_signed(4, 5),
    7 => to_signed(4, 5),
    8 => to_signed(4, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(4, 5),
    12 => to_signed(4, 5),
    13 => to_signed(4, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-2, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-3, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-4, 5),
    59 => to_signed(-4, 5),
    60 => to_signed(-5, 5),
    61 => to_signed(-5, 5),
    62 => to_signed(-5, 5),
    63 => to_signed(-6, 5)
  );

  constant LUT_0_10_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_11_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(0, 5),
    54 => to_signed(0, 5),
    55 => to_signed(0, 5),
    56 => to_signed(0, 5),
    57 => to_signed(0, 5),
    58 => to_signed(0, 5),
    59 => to_signed(0, 5),
    60 => to_signed(1, 5),
    61 => to_signed(1, 5),
    62 => to_signed(1, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_11_1_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-4, 5),
    44 => to_signed(-4, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-5, 5),
    47 => to_signed(-5, 5),
    48 => to_signed(-5, 5),
    49 => to_signed(-6, 5),
    50 => to_signed(-6, 5),
    51 => to_signed(-7, 5),
    52 => to_signed(-7, 5),
    53 => to_signed(-7, 5),
    54 => to_signed(-8, 5),
    55 => to_signed(-8, 5),
    56 => to_signed(-9, 5),
    57 => to_signed(-9, 5),
    58 => to_signed(-9, 5),
    59 => to_signed(-10, 5),
    60 => to_signed(-10, 5),
    61 => to_signed(-11, 5),
    62 => to_signed(-11, 5),
    63 => to_signed(-11, 5)
  );

  constant LUT_0_11_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(3, 5),
    9 => to_signed(3, 5),
    10 => to_signed(3, 5),
    11 => to_signed(3, 5),
    12 => to_signed(3, 5),
    13 => to_signed(3, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-4, 5),
    59 => to_signed(-4, 5),
    60 => to_signed(-4, 5),
    61 => to_signed(-4, 5),
    62 => to_signed(-4, 5),
    63 => to_signed(-4, 5)
  );

  constant LUT_0_11_3_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(3, 5),
    5 => to_signed(3, 5),
    6 => to_signed(3, 5),
    7 => to_signed(4, 5),
    8 => to_signed(4, 5),
    9 => to_signed(4, 5),
    10 => to_signed(5, 5),
    11 => to_signed(5, 5),
    12 => to_signed(5, 5),
    13 => to_signed(5, 5),
    14 => to_signed(5, 5),
    15 => to_signed(5, 5),
    16 => to_signed(4, 5),
    17 => to_signed(4, 5),
    18 => to_signed(4, 5),
    19 => to_signed(3, 5),
    20 => to_signed(3, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-2, 5),
    33 => to_signed(-2, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-3, 5),
    37 => to_signed(-3, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-3, 5),
    43 => to_signed(-3, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-4, 5),
    46 => to_signed(-4, 5),
    47 => to_signed(-4, 5),
    48 => to_signed(-4, 5),
    49 => to_signed(-4, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-3, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_11_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(4, 5),
    58 => to_signed(4, 5),
    59 => to_signed(4, 5),
    60 => to_signed(4, 5),
    61 => to_signed(5, 5),
    62 => to_signed(5, 5),
    63 => to_signed(5, 5)
  );

  constant LUT_0_11_5_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-3, 5),
    57 => to_signed(-3, 5),
    58 => to_signed(-3, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-4, 5),
    63 => to_signed(-4, 5)
  );

  constant LUT_0_11_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_11_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-3, 5),
    9 => to_signed(-3, 5),
    10 => to_signed(-3, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-3, 5),
    13 => to_signed(-3, 5),
    14 => to_signed(-3, 5),
    15 => to_signed(-3, 5),
    16 => to_signed(-3, 5),
    17 => to_signed(-3, 5),
    18 => to_signed(-3, 5),
    19 => to_signed(-3, 5),
    20 => to_signed(-3, 5),
    21 => to_signed(-3, 5),
    22 => to_signed(-3, 5),
    23 => to_signed(-3, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-2, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(1, 5),
    34 => to_signed(1, 5),
    35 => to_signed(2, 5),
    36 => to_signed(2, 5),
    37 => to_signed(2, 5),
    38 => to_signed(3, 5),
    39 => to_signed(3, 5),
    40 => to_signed(4, 5),
    41 => to_signed(4, 5),
    42 => to_signed(5, 5),
    43 => to_signed(5, 5),
    44 => to_signed(6, 5),
    45 => to_signed(6, 5),
    46 => to_signed(6, 5),
    47 => to_signed(7, 5),
    48 => to_signed(7, 5),
    49 => to_signed(8, 5),
    50 => to_signed(8, 5),
    51 => to_signed(8, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(10, 5),
    57 => to_signed(11, 5),
    58 => to_signed(11, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(13, 5),
    62 => to_signed(13, 5),
    63 => to_signed(13, 5)
  );

  constant LUT_0_12_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-3, 5),
    57 => to_signed(-3, 5),
    58 => to_signed(-3, 5),
    59 => to_signed(-4, 5),
    60 => to_signed(-4, 5),
    61 => to_signed(-4, 5),
    62 => to_signed(-4, 5),
    63 => to_signed(-4, 5)
  );

  constant LUT_0_12_1_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(2, 5),
    46 => to_signed(2, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(3, 5),
    53 => to_signed(3, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_12_2_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-1, 5),
    48 => to_signed(-1, 5),
    49 => to_signed(-1, 5),
    50 => to_signed(-1, 5),
    51 => to_signed(-1, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_12_3_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_12_4_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(2, 5),
    55 => to_signed(2, 5),
    56 => to_signed(2, 5),
    57 => to_signed(2, 5),
    58 => to_signed(2, 5),
    59 => to_signed(3, 5),
    60 => to_signed(3, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_12_5_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(-1, 5),
    17 => to_signed(-1, 5),
    18 => to_signed(-1, 5),
    19 => to_signed(-1, 5),
    20 => to_signed(-1, 5),
    21 => to_signed(-1, 5),
    22 => to_signed(-1, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(1, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(2, 5),
    43 => to_signed(3, 5),
    44 => to_signed(3, 5),
    45 => to_signed(3, 5),
    46 => to_signed(3, 5),
    47 => to_signed(4, 5),
    48 => to_signed(4, 5),
    49 => to_signed(4, 5),
    50 => to_signed(5, 5),
    51 => to_signed(5, 5),
    52 => to_signed(5, 5),
    53 => to_signed(5, 5),
    54 => to_signed(6, 5),
    55 => to_signed(6, 5),
    56 => to_signed(6, 5),
    57 => to_signed(7, 5),
    58 => to_signed(7, 5),
    59 => to_signed(7, 5),
    60 => to_signed(8, 5),
    61 => to_signed(8, 5),
    62 => to_signed(8, 5),
    63 => to_signed(9, 5)
  );

  constant LUT_0_12_6_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-2, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-3, 5),
    45 => to_signed(-3, 5),
    46 => to_signed(-3, 5),
    47 => to_signed(-3, 5),
    48 => to_signed(-3, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-4, 5),
    51 => to_signed(-4, 5),
    52 => to_signed(-4, 5),
    53 => to_signed(-4, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-5, 5),
    57 => to_signed(-5, 5),
    58 => to_signed(-5, 5),
    59 => to_signed(-5, 5),
    60 => to_signed(-6, 5),
    61 => to_signed(-6, 5),
    62 => to_signed(-6, 5),
    63 => to_signed(-6, 5)
  );

  constant LUT_0_12_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(2, 5),
    17 => to_signed(2, 5),
    18 => to_signed(2, 5),
    19 => to_signed(2, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(2, 5),
    25 => to_signed(2, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-2, 5),
    39 => to_signed(-2, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-3, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-4, 5),
    44 => to_signed(-5, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-6, 5),
    47 => to_signed(-6, 5),
    48 => to_signed(-7, 5),
    49 => to_signed(-7, 5),
    50 => to_signed(-8, 5),
    51 => to_signed(-8, 5),
    52 => to_signed(-9, 5),
    53 => to_signed(-9, 5),
    54 => to_signed(-10, 5),
    55 => to_signed(-10, 5),
    56 => to_signed(-11, 5),
    57 => to_signed(-11, 5),
    58 => to_signed(-12, 5),
    59 => to_signed(-12, 5),
    60 => to_signed(-13, 5),
    61 => to_signed(-13, 5),
    62 => to_signed(-14, 5),
    63 => to_signed(-14, 5)
  );

  constant LUT_0_13_0_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(0, 5),
    53 => to_signed(0, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-1, 5),
    61 => to_signed(-1, 5),
    62 => to_signed(-1, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_13_1_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-2, 5),
    43 => to_signed(-2, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-3, 5),
    59 => to_signed(-3, 5),
    60 => to_signed(-3, 5),
    61 => to_signed(-3, 5),
    62 => to_signed(-3, 5),
    63 => to_signed(-3, 5)
  );

  constant LUT_0_13_2_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(0, 5),
    43 => to_signed(0, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(1, 5),
    57 => to_signed(1, 5),
    58 => to_signed(1, 5),
    59 => to_signed(1, 5),
    60 => to_signed(1, 5),
    61 => to_signed(0, 5),
    62 => to_signed(0, 5),
    63 => to_signed(0, 5)
  );

  constant LUT_0_13_3_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(0, 5),
    11 => to_signed(0, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(1, 5),
    40 => to_signed(1, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(2, 5),
    48 => to_signed(2, 5),
    49 => to_signed(2, 5),
    50 => to_signed(2, 5),
    51 => to_signed(2, 5),
    52 => to_signed(2, 5),
    53 => to_signed(2, 5),
    54 => to_signed(3, 5),
    55 => to_signed(3, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(3, 5),
    59 => to_signed(3, 5),
    60 => to_signed(4, 5),
    61 => to_signed(4, 5),
    62 => to_signed(4, 5),
    63 => to_signed(4, 5)
  );

  constant LUT_0_13_4_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(1, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-2, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-3, 5),
    55 => to_signed(-3, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-4, 5),
    58 => to_signed(-4, 5),
    59 => to_signed(-4, 5),
    60 => to_signed(-5, 5),
    61 => to_signed(-5, 5),
    62 => to_signed(-5, 5),
    63 => to_signed(-5, 5)
  );

  constant LUT_0_13_5_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(1, 5),
    2 => to_signed(1, 5),
    3 => to_signed(2, 5),
    4 => to_signed(2, 5),
    5 => to_signed(2, 5),
    6 => to_signed(2, 5),
    7 => to_signed(2, 5),
    8 => to_signed(2, 5),
    9 => to_signed(2, 5),
    10 => to_signed(2, 5),
    11 => to_signed(2, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(2, 5),
    15 => to_signed(2, 5),
    16 => to_signed(2, 5),
    17 => to_signed(1, 5),
    18 => to_signed(1, 5),
    19 => to_signed(1, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(-1, 5),
    39 => to_signed(-1, 5),
    40 => to_signed(-1, 5),
    41 => to_signed(-1, 5),
    42 => to_signed(-1, 5),
    43 => to_signed(-1, 5),
    44 => to_signed(-1, 5),
    45 => to_signed(-2, 5),
    46 => to_signed(-2, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(-2, 5),
    53 => to_signed(-2, 5),
    54 => to_signed(-2, 5),
    55 => to_signed(-2, 5),
    56 => to_signed(-2, 5),
    57 => to_signed(-2, 5),
    58 => to_signed(-2, 5),
    59 => to_signed(-2, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_13_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(0, 5),
    5 => to_signed(0, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(0, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(0, 5),
    13 => to_signed(0, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(0, 5),
    24 => to_signed(0, 5),
    25 => to_signed(0, 5),
    26 => to_signed(0, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(1, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(1, 5),
    45 => to_signed(1, 5),
    46 => to_signed(1, 5),
    47 => to_signed(1, 5),
    48 => to_signed(1, 5),
    49 => to_signed(1, 5),
    50 => to_signed(1, 5),
    51 => to_signed(1, 5),
    52 => to_signed(1, 5),
    53 => to_signed(1, 5),
    54 => to_signed(1, 5),
    55 => to_signed(1, 5),
    56 => to_signed(1, 5),
    57 => to_signed(1, 5),
    58 => to_signed(1, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(2, 5),
    62 => to_signed(2, 5),
    63 => to_signed(2, 5)
  );

  constant LUT_0_13_7_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(0, 5),
    2 => to_signed(0, 5),
    3 => to_signed(0, 5),
    4 => to_signed(1, 5),
    5 => to_signed(1, 5),
    6 => to_signed(1, 5),
    7 => to_signed(1, 5),
    8 => to_signed(1, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(1, 5),
    13 => to_signed(1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(1, 5),
    16 => to_signed(1, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(0, 5),
    34 => to_signed(0, 5),
    35 => to_signed(0, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(0, 5),
    39 => to_signed(0, 5),
    40 => to_signed(0, 5),
    41 => to_signed(0, 5),
    42 => to_signed(1, 5),
    43 => to_signed(1, 5),
    44 => to_signed(0, 5),
    45 => to_signed(0, 5),
    46 => to_signed(0, 5),
    47 => to_signed(0, 5),
    48 => to_signed(0, 5),
    49 => to_signed(0, 5),
    50 => to_signed(0, 5),
    51 => to_signed(0, 5),
    52 => to_signed(-1, 5),
    53 => to_signed(-1, 5),
    54 => to_signed(-1, 5),
    55 => to_signed(-1, 5),
    56 => to_signed(-1, 5),
    57 => to_signed(-1, 5),
    58 => to_signed(-1, 5),
    59 => to_signed(-1, 5),
    60 => to_signed(-2, 5),
    61 => to_signed(-2, 5),
    62 => to_signed(-2, 5),
    63 => to_signed(-2, 5)
  );

  constant LUT_0_14_0_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-2, 5),
    9 => to_signed(-2, 5),
    10 => to_signed(-2, 5),
    11 => to_signed(-2, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(1, 5),
    21 => to_signed(1, 5),
    22 => to_signed(1, 5),
    23 => to_signed(1, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(-2, 5),
    32 => to_signed(-2, 5),
    33 => to_signed(-2, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-1, 5),
    37 => to_signed(-1, 5),
    38 => to_signed(0, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(2, 5),
    42 => to_signed(3, 5),
    43 => to_signed(4, 5),
    44 => to_signed(5, 5),
    45 => to_signed(5, 5),
    46 => to_signed(6, 5),
    47 => to_signed(7, 5),
    48 => to_signed(7, 5),
    49 => to_signed(8, 5),
    50 => to_signed(8, 5),
    51 => to_signed(9, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(11, 5),
    57 => to_signed(11, 5),
    58 => to_signed(12, 5),
    59 => to_signed(12, 5),
    60 => to_signed(13, 5),
    61 => to_signed(14, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_14_1_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-2, 5),
    7 => to_signed(-2, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(0, 5),
    15 => to_signed(0, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(0, 5),
    19 => to_signed(0, 5),
    20 => to_signed(0, 5),
    21 => to_signed(0, 5),
    22 => to_signed(0, 5),
    23 => to_signed(-1, 5),
    24 => to_signed(-1, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-2, 5),
    32 => to_signed(-2, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(0, 5),
    37 => to_signed(0, 5),
    38 => to_signed(1, 5),
    39 => to_signed(1, 5),
    40 => to_signed(2, 5),
    41 => to_signed(3, 5),
    42 => to_signed(3, 5),
    43 => to_signed(4, 5),
    44 => to_signed(4, 5),
    45 => to_signed(5, 5),
    46 => to_signed(5, 5),
    47 => to_signed(5, 5),
    48 => to_signed(5, 5),
    49 => to_signed(5, 5),
    50 => to_signed(5, 5),
    51 => to_signed(5, 5),
    52 => to_signed(5, 5),
    53 => to_signed(4, 5),
    54 => to_signed(4, 5),
    55 => to_signed(4, 5),
    56 => to_signed(3, 5),
    57 => to_signed(3, 5),
    58 => to_signed(2, 5),
    59 => to_signed(2, 5),
    60 => to_signed(2, 5),
    61 => to_signed(3, 5),
    62 => to_signed(3, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_14_2_DATA : lut_array_t_0 := (
    0 => to_signed(-4, 5),
    1 => to_signed(-4, 5),
    2 => to_signed(-5, 5),
    3 => to_signed(-5, 5),
    4 => to_signed(-5, 5),
    5 => to_signed(-5, 5),
    6 => to_signed(-5, 5),
    7 => to_signed(-5, 5),
    8 => to_signed(-6, 5),
    9 => to_signed(-6, 5),
    10 => to_signed(-6, 5),
    11 => to_signed(-6, 5),
    12 => to_signed(-6, 5),
    13 => to_signed(-7, 5),
    14 => to_signed(-7, 5),
    15 => to_signed(-8, 5),
    16 => to_signed(-9, 5),
    17 => to_signed(-9, 5),
    18 => to_signed(-9, 5),
    19 => to_signed(-9, 5),
    20 => to_signed(-9, 5),
    21 => to_signed(-9, 5),
    22 => to_signed(-9, 5),
    23 => to_signed(-8, 5),
    24 => to_signed(-8, 5),
    25 => to_signed(-7, 5),
    26 => to_signed(-6, 5),
    27 => to_signed(-5, 5),
    28 => to_signed(-4, 5),
    29 => to_signed(-3, 5),
    30 => to_signed(-2, 5),
    31 => to_signed(-1, 5),
    32 => to_signed(1, 5),
    33 => to_signed(2, 5),
    34 => to_signed(3, 5),
    35 => to_signed(4, 5),
    36 => to_signed(6, 5),
    37 => to_signed(7, 5),
    38 => to_signed(7, 5),
    39 => to_signed(8, 5),
    40 => to_signed(8, 5),
    41 => to_signed(8, 5),
    42 => to_signed(8, 5),
    43 => to_signed(8, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(7, 5),
    47 => to_signed(7, 5),
    48 => to_signed(7, 5),
    49 => to_signed(8, 5),
    50 => to_signed(8, 5),
    51 => to_signed(8, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(9, 5),
    55 => to_signed(9, 5),
    56 => to_signed(10, 5),
    57 => to_signed(10, 5),
    58 => to_signed(11, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(13, 5),
    62 => to_signed(14, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_14_3_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(0, 5),
    7 => to_signed(0, 5),
    8 => to_signed(0, 5),
    9 => to_signed(1, 5),
    10 => to_signed(1, 5),
    11 => to_signed(1, 5),
    12 => to_signed(2, 5),
    13 => to_signed(2, 5),
    14 => to_signed(3, 5),
    15 => to_signed(3, 5),
    16 => to_signed(3, 5),
    17 => to_signed(4, 5),
    18 => to_signed(4, 5),
    19 => to_signed(5, 5),
    20 => to_signed(6, 5),
    21 => to_signed(6, 5),
    22 => to_signed(7, 5),
    23 => to_signed(7, 5),
    24 => to_signed(8, 5),
    25 => to_signed(8, 5),
    26 => to_signed(8, 5),
    27 => to_signed(8, 5),
    28 => to_signed(7, 5),
    29 => to_signed(7, 5),
    30 => to_signed(6, 5),
    31 => to_signed(4, 5),
    32 => to_signed(3, 5),
    33 => to_signed(1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-4, 5),
    37 => to_signed(-5, 5),
    38 => to_signed(-7, 5),
    39 => to_signed(-7, 5),
    40 => to_signed(-8, 5),
    41 => to_signed(-8, 5),
    42 => to_signed(-7, 5),
    43 => to_signed(-7, 5),
    44 => to_signed(-6, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-5, 5),
    47 => to_signed(-4, 5),
    48 => to_signed(-4, 5),
    49 => to_signed(-3, 5),
    50 => to_signed(-2, 5),
    51 => to_signed(-2, 5),
    52 => to_signed(0, 5),
    53 => to_signed(1, 5),
    54 => to_signed(2, 5),
    55 => to_signed(4, 5),
    56 => to_signed(5, 5),
    57 => to_signed(6, 5),
    58 => to_signed(7, 5),
    59 => to_signed(7, 5),
    60 => to_signed(6, 5),
    61 => to_signed(5, 5),
    62 => to_signed(4, 5),
    63 => to_signed(3, 5)
  );

  constant LUT_0_14_4_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-3, 5),
    2 => to_signed(-3, 5),
    3 => to_signed(-3, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-3, 5),
    8 => to_signed(-3, 5),
    9 => to_signed(-3, 5),
    10 => to_signed(-3, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-2, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-1, 5),
    16 => to_signed(0, 5),
    17 => to_signed(0, 5),
    18 => to_signed(1, 5),
    19 => to_signed(2, 5),
    20 => to_signed(3, 5),
    21 => to_signed(4, 5),
    22 => to_signed(5, 5),
    23 => to_signed(6, 5),
    24 => to_signed(7, 5),
    25 => to_signed(7, 5),
    26 => to_signed(7, 5),
    27 => to_signed(7, 5),
    28 => to_signed(6, 5),
    29 => to_signed(5, 5),
    30 => to_signed(4, 5),
    31 => to_signed(3, 5),
    32 => to_signed(1, 5),
    33 => to_signed(0, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-3, 5),
    36 => to_signed(-4, 5),
    37 => to_signed(-5, 5),
    38 => to_signed(-5, 5),
    39 => to_signed(-5, 5),
    40 => to_signed(-4, 5),
    41 => to_signed(-2, 5),
    42 => to_signed(0, 5),
    43 => to_signed(2, 5),
    44 => to_signed(4, 5),
    45 => to_signed(7, 5),
    46 => to_signed(9, 5),
    47 => to_signed(12, 5),
    48 => to_signed(14, 5),
    49 => to_signed(15, 5),
    50 => to_signed(15, 5),
    51 => to_signed(15, 5),
    52 => to_signed(15, 5),
    53 => to_signed(15, 5),
    54 => to_signed(15, 5),
    55 => to_signed(15, 5),
    56 => to_signed(15, 5),
    57 => to_signed(15, 5),
    58 => to_signed(14, 5),
    59 => to_signed(13, 5),
    60 => to_signed(12, 5),
    61 => to_signed(11, 5),
    62 => to_signed(11, 5),
    63 => to_signed(10, 5)
  );

  constant LUT_0_14_5_DATA : lut_array_t_0 := (
    0 => to_signed(7, 5),
    1 => to_signed(8, 5),
    2 => to_signed(9, 5),
    3 => to_signed(10, 5),
    4 => to_signed(11, 5),
    5 => to_signed(11, 5),
    6 => to_signed(12, 5),
    7 => to_signed(12, 5),
    8 => to_signed(12, 5),
    9 => to_signed(12, 5),
    10 => to_signed(12, 5),
    11 => to_signed(12, 5),
    12 => to_signed(11, 5),
    13 => to_signed(11, 5),
    14 => to_signed(10, 5),
    15 => to_signed(10, 5),
    16 => to_signed(9, 5),
    17 => to_signed(8, 5),
    18 => to_signed(8, 5),
    19 => to_signed(7, 5),
    20 => to_signed(7, 5),
    21 => to_signed(7, 5),
    22 => to_signed(7, 5),
    23 => to_signed(7, 5),
    24 => to_signed(7, 5),
    25 => to_signed(6, 5),
    26 => to_signed(6, 5),
    27 => to_signed(5, 5),
    28 => to_signed(4, 5),
    29 => to_signed(3, 5),
    30 => to_signed(2, 5),
    31 => to_signed(1, 5),
    32 => to_signed(0, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-3, 5),
    35 => to_signed(-4, 5),
    36 => to_signed(-5, 5),
    37 => to_signed(-6, 5),
    38 => to_signed(-7, 5),
    39 => to_signed(-8, 5),
    40 => to_signed(-8, 5),
    41 => to_signed(-9, 5),
    42 => to_signed(-9, 5),
    43 => to_signed(-10, 5),
    44 => to_signed(-11, 5),
    45 => to_signed(-12, 5),
    46 => to_signed(-13, 5),
    47 => to_signed(-14, 5),
    48 => to_signed(-15, 5),
    49 => to_signed(-16, 5),
    50 => to_signed(-16, 5),
    51 => to_signed(-16, 5),
    52 => to_signed(-16, 5),
    53 => to_signed(-16, 5),
    54 => to_signed(-16, 5),
    55 => to_signed(-16, 5),
    56 => to_signed(-16, 5),
    57 => to_signed(-16, 5),
    58 => to_signed(-16, 5),
    59 => to_signed(-16, 5),
    60 => to_signed(-16, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_14_6_DATA : lut_array_t_0 := (
    0 => to_signed(0, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-4, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-3, 5),
    12 => to_signed(-2, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(1, 5),
    15 => to_signed(3, 5),
    16 => to_signed(5, 5),
    17 => to_signed(8, 5),
    18 => to_signed(10, 5),
    19 => to_signed(12, 5),
    20 => to_signed(14, 5),
    21 => to_signed(15, 5),
    22 => to_signed(15, 5),
    23 => to_signed(15, 5),
    24 => to_signed(15, 5),
    25 => to_signed(15, 5),
    26 => to_signed(15, 5),
    27 => to_signed(15, 5),
    28 => to_signed(14, 5),
    29 => to_signed(13, 5),
    30 => to_signed(11, 5),
    31 => to_signed(8, 5),
    32 => to_signed(6, 5),
    33 => to_signed(4, 5),
    34 => to_signed(2, 5),
    35 => to_signed(-1, 5),
    36 => to_signed(-3, 5),
    37 => to_signed(-4, 5),
    38 => to_signed(-6, 5),
    39 => to_signed(-8, 5),
    40 => to_signed(-9, 5),
    41 => to_signed(-10, 5),
    42 => to_signed(-11, 5),
    43 => to_signed(-11, 5),
    44 => to_signed(-12, 5),
    45 => to_signed(-13, 5),
    46 => to_signed(-13, 5),
    47 => to_signed(-14, 5),
    48 => to_signed(-15, 5),
    49 => to_signed(-16, 5),
    50 => to_signed(-16, 5),
    51 => to_signed(-16, 5),
    52 => to_signed(-16, 5),
    53 => to_signed(-16, 5),
    54 => to_signed(-16, 5),
    55 => to_signed(-16, 5),
    56 => to_signed(-16, 5),
    57 => to_signed(-16, 5),
    58 => to_signed(-16, 5),
    59 => to_signed(-16, 5),
    60 => to_signed(-16, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  constant LUT_0_14_7_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-3, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-4, 5),
    12 => to_signed(-5, 5),
    13 => to_signed(-6, 5),
    14 => to_signed(-6, 5),
    15 => to_signed(-7, 5),
    16 => to_signed(-8, 5),
    17 => to_signed(-8, 5),
    18 => to_signed(-9, 5),
    19 => to_signed(-9, 5),
    20 => to_signed(-9, 5),
    21 => to_signed(-9, 5),
    22 => to_signed(-8, 5),
    23 => to_signed(-7, 5),
    24 => to_signed(-6, 5),
    25 => to_signed(-4, 5),
    26 => to_signed(-3, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(0, 5),
    29 => to_signed(2, 5),
    30 => to_signed(3, 5),
    31 => to_signed(4, 5),
    32 => to_signed(5, 5),
    33 => to_signed(6, 5),
    34 => to_signed(6, 5),
    35 => to_signed(6, 5),
    36 => to_signed(6, 5),
    37 => to_signed(6, 5),
    38 => to_signed(5, 5),
    39 => to_signed(4, 5),
    40 => to_signed(3, 5),
    41 => to_signed(3, 5),
    42 => to_signed(2, 5),
    43 => to_signed(1, 5),
    44 => to_signed(0, 5),
    45 => to_signed(-1, 5),
    46 => to_signed(-1, 5),
    47 => to_signed(-2, 5),
    48 => to_signed(-2, 5),
    49 => to_signed(-2, 5),
    50 => to_signed(-3, 5),
    51 => to_signed(-3, 5),
    52 => to_signed(-3, 5),
    53 => to_signed(-3, 5),
    54 => to_signed(-4, 5),
    55 => to_signed(-4, 5),
    56 => to_signed(-4, 5),
    57 => to_signed(-5, 5),
    58 => to_signed(-6, 5),
    59 => to_signed(-7, 5),
    60 => to_signed(-8, 5),
    61 => to_signed(-9, 5),
    62 => to_signed(-10, 5),
    63 => to_signed(-11, 5)
  );

  constant LUT_0_15_0_DATA : lut_array_t_0 := (
    0 => to_signed(-3, 5),
    1 => to_signed(-3, 5),
    2 => to_signed(-4, 5),
    3 => to_signed(-5, 5),
    4 => to_signed(-6, 5),
    5 => to_signed(-7, 5),
    6 => to_signed(-7, 5),
    7 => to_signed(-8, 5),
    8 => to_signed(-9, 5),
    9 => to_signed(-9, 5),
    10 => to_signed(-10, 5),
    11 => to_signed(-10, 5),
    12 => to_signed(-11, 5),
    13 => to_signed(-11, 5),
    14 => to_signed(-11, 5),
    15 => to_signed(-11, 5),
    16 => to_signed(-11, 5),
    17 => to_signed(-10, 5),
    18 => to_signed(-10, 5),
    19 => to_signed(-9, 5),
    20 => to_signed(-8, 5),
    21 => to_signed(-7, 5),
    22 => to_signed(-6, 5),
    23 => to_signed(-5, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(1, 5),
    29 => to_signed(1, 5),
    30 => to_signed(2, 5),
    31 => to_signed(3, 5),
    32 => to_signed(3, 5),
    33 => to_signed(3, 5),
    34 => to_signed(4, 5),
    35 => to_signed(4, 5),
    36 => to_signed(4, 5),
    37 => to_signed(4, 5),
    38 => to_signed(4, 5),
    39 => to_signed(5, 5),
    40 => to_signed(5, 5),
    41 => to_signed(5, 5),
    42 => to_signed(6, 5),
    43 => to_signed(6, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(8, 5),
    47 => to_signed(8, 5),
    48 => to_signed(9, 5),
    49 => to_signed(9, 5),
    50 => to_signed(9, 5),
    51 => to_signed(10, 5),
    52 => to_signed(10, 5),
    53 => to_signed(11, 5),
    54 => to_signed(11, 5),
    55 => to_signed(11, 5),
    56 => to_signed(12, 5),
    57 => to_signed(12, 5),
    58 => to_signed(12, 5),
    59 => to_signed(12, 5),
    60 => to_signed(12, 5),
    61 => to_signed(12, 5),
    62 => to_signed(12, 5),
    63 => to_signed(12, 5)
  );

  constant LUT_0_15_1_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-1, 5),
    3 => to_signed(-1, 5),
    4 => to_signed(-1, 5),
    5 => to_signed(-1, 5),
    6 => to_signed(-1, 5),
    7 => to_signed(-1, 5),
    8 => to_signed(-1, 5),
    9 => to_signed(-1, 5),
    10 => to_signed(-1, 5),
    11 => to_signed(-1, 5),
    12 => to_signed(-1, 5),
    13 => to_signed(-1, 5),
    14 => to_signed(-1, 5),
    15 => to_signed(-2, 5),
    16 => to_signed(-2, 5),
    17 => to_signed(-2, 5),
    18 => to_signed(-2, 5),
    19 => to_signed(-2, 5),
    20 => to_signed(-2, 5),
    21 => to_signed(-2, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-2, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(-1, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(0, 5),
    34 => to_signed(1, 5),
    35 => to_signed(1, 5),
    36 => to_signed(1, 5),
    37 => to_signed(2, 5),
    38 => to_signed(2, 5),
    39 => to_signed(3, 5),
    40 => to_signed(3, 5),
    41 => to_signed(3, 5),
    42 => to_signed(4, 5),
    43 => to_signed(4, 5),
    44 => to_signed(5, 5),
    45 => to_signed(5, 5),
    46 => to_signed(6, 5),
    47 => to_signed(6, 5),
    48 => to_signed(7, 5),
    49 => to_signed(7, 5),
    50 => to_signed(8, 5),
    51 => to_signed(8, 5),
    52 => to_signed(9, 5),
    53 => to_signed(9, 5),
    54 => to_signed(10, 5),
    55 => to_signed(10, 5),
    56 => to_signed(11, 5),
    57 => to_signed(12, 5),
    58 => to_signed(12, 5),
    59 => to_signed(13, 5),
    60 => to_signed(13, 5),
    61 => to_signed(14, 5),
    62 => to_signed(14, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_15_2_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-3, 5),
    3 => to_signed(-3, 5),
    4 => to_signed(-4, 5),
    5 => to_signed(-4, 5),
    6 => to_signed(-5, 5),
    7 => to_signed(-5, 5),
    8 => to_signed(-6, 5),
    9 => to_signed(-6, 5),
    10 => to_signed(-6, 5),
    11 => to_signed(-7, 5),
    12 => to_signed(-7, 5),
    13 => to_signed(-7, 5),
    14 => to_signed(-7, 5),
    15 => to_signed(-7, 5),
    16 => to_signed(-6, 5),
    17 => to_signed(-6, 5),
    18 => to_signed(-6, 5),
    19 => to_signed(-5, 5),
    20 => to_signed(-5, 5),
    21 => to_signed(-4, 5),
    22 => to_signed(-4, 5),
    23 => to_signed(-4, 5),
    24 => to_signed(-3, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-2, 5),
    27 => to_signed(-1, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(1, 5),
    32 => to_signed(2, 5),
    33 => to_signed(2, 5),
    34 => to_signed(3, 5),
    35 => to_signed(3, 5),
    36 => to_signed(4, 5),
    37 => to_signed(4, 5),
    38 => to_signed(5, 5),
    39 => to_signed(5, 5),
    40 => to_signed(6, 5),
    41 => to_signed(6, 5),
    42 => to_signed(6, 5),
    43 => to_signed(7, 5),
    44 => to_signed(7, 5),
    45 => to_signed(7, 5),
    46 => to_signed(8, 5),
    47 => to_signed(8, 5),
    48 => to_signed(8, 5),
    49 => to_signed(8, 5),
    50 => to_signed(9, 5),
    51 => to_signed(9, 5),
    52 => to_signed(9, 5),
    53 => to_signed(10, 5),
    54 => to_signed(10, 5),
    55 => to_signed(11, 5),
    56 => to_signed(11, 5),
    57 => to_signed(12, 5),
    58 => to_signed(12, 5),
    59 => to_signed(13, 5),
    60 => to_signed(13, 5),
    61 => to_signed(14, 5),
    62 => to_signed(14, 5),
    63 => to_signed(14, 5)
  );

  constant LUT_0_15_3_DATA : lut_array_t_0 := (
    0 => to_signed(-4, 5),
    1 => to_signed(-5, 5),
    2 => to_signed(-6, 5),
    3 => to_signed(-7, 5),
    4 => to_signed(-9, 5),
    5 => to_signed(-10, 5),
    6 => to_signed(-11, 5),
    7 => to_signed(-12, 5),
    8 => to_signed(-13, 5),
    9 => to_signed(-14, 5),
    10 => to_signed(-14, 5),
    11 => to_signed(-15, 5),
    12 => to_signed(-15, 5),
    13 => to_signed(-14, 5),
    14 => to_signed(-14, 5),
    15 => to_signed(-13, 5),
    16 => to_signed(-13, 5),
    17 => to_signed(-12, 5),
    18 => to_signed(-11, 5),
    19 => to_signed(-10, 5),
    20 => to_signed(-9, 5),
    21 => to_signed(-7, 5),
    22 => to_signed(-6, 5),
    23 => to_signed(-5, 5),
    24 => to_signed(-4, 5),
    25 => to_signed(-3, 5),
    26 => to_signed(-3, 5),
    27 => to_signed(-2, 5),
    28 => to_signed(-1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(2, 5),
    33 => to_signed(3, 5),
    34 => to_signed(3, 5),
    35 => to_signed(4, 5),
    36 => to_signed(4, 5),
    37 => to_signed(5, 5),
    38 => to_signed(6, 5),
    39 => to_signed(6, 5),
    40 => to_signed(7, 5),
    41 => to_signed(8, 5),
    42 => to_signed(8, 5),
    43 => to_signed(9, 5),
    44 => to_signed(10, 5),
    45 => to_signed(10, 5),
    46 => to_signed(11, 5),
    47 => to_signed(12, 5),
    48 => to_signed(12, 5),
    49 => to_signed(13, 5),
    50 => to_signed(13, 5),
    51 => to_signed(14, 5),
    52 => to_signed(15, 5),
    53 => to_signed(15, 5),
    54 => to_signed(15, 5),
    55 => to_signed(15, 5),
    56 => to_signed(15, 5),
    57 => to_signed(15, 5),
    58 => to_signed(15, 5),
    59 => to_signed(15, 5),
    60 => to_signed(15, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_15_4_DATA : lut_array_t_0 := (
    0 => to_signed(-1, 5),
    1 => to_signed(-1, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-2, 5),
    5 => to_signed(-2, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-3, 5),
    8 => to_signed(-3, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-4, 5),
    11 => to_signed(-4, 5),
    12 => to_signed(-5, 5),
    13 => to_signed(-5, 5),
    14 => to_signed(-6, 5),
    15 => to_signed(-6, 5),
    16 => to_signed(-7, 5),
    17 => to_signed(-7, 5),
    18 => to_signed(-7, 5),
    19 => to_signed(-8, 5),
    20 => to_signed(-7, 5),
    21 => to_signed(-7, 5),
    22 => to_signed(-7, 5),
    23 => to_signed(-6, 5),
    24 => to_signed(-6, 5),
    25 => to_signed(-5, 5),
    26 => to_signed(-5, 5),
    27 => to_signed(-4, 5),
    28 => to_signed(-3, 5),
    29 => to_signed(-2, 5),
    30 => to_signed(-1, 5),
    31 => to_signed(0, 5),
    32 => to_signed(1, 5),
    33 => to_signed(1, 5),
    34 => to_signed(2, 5),
    35 => to_signed(3, 5),
    36 => to_signed(4, 5),
    37 => to_signed(5, 5),
    38 => to_signed(6, 5),
    39 => to_signed(7, 5),
    40 => to_signed(8, 5),
    41 => to_signed(9, 5),
    42 => to_signed(9, 5),
    43 => to_signed(10, 5),
    44 => to_signed(11, 5),
    45 => to_signed(12, 5),
    46 => to_signed(12, 5),
    47 => to_signed(13, 5),
    48 => to_signed(13, 5),
    49 => to_signed(14, 5),
    50 => to_signed(14, 5),
    51 => to_signed(15, 5),
    52 => to_signed(15, 5),
    53 => to_signed(15, 5),
    54 => to_signed(15, 5),
    55 => to_signed(14, 5),
    56 => to_signed(14, 5),
    57 => to_signed(14, 5),
    58 => to_signed(14, 5),
    59 => to_signed(14, 5),
    60 => to_signed(14, 5),
    61 => to_signed(15, 5),
    62 => to_signed(15, 5),
    63 => to_signed(15, 5)
  );

  constant LUT_0_15_5_DATA : lut_array_t_0 := (
    0 => to_signed(1, 5),
    1 => to_signed(2, 5),
    2 => to_signed(2, 5),
    3 => to_signed(2, 5),
    4 => to_signed(3, 5),
    5 => to_signed(3, 5),
    6 => to_signed(3, 5),
    7 => to_signed(3, 5),
    8 => to_signed(3, 5),
    9 => to_signed(4, 5),
    10 => to_signed(4, 5),
    11 => to_signed(4, 5),
    12 => to_signed(4, 5),
    13 => to_signed(4, 5),
    14 => to_signed(4, 5),
    15 => to_signed(4, 5),
    16 => to_signed(3, 5),
    17 => to_signed(3, 5),
    18 => to_signed(3, 5),
    19 => to_signed(3, 5),
    20 => to_signed(2, 5),
    21 => to_signed(2, 5),
    22 => to_signed(2, 5),
    23 => to_signed(2, 5),
    24 => to_signed(1, 5),
    25 => to_signed(1, 5),
    26 => to_signed(1, 5),
    27 => to_signed(1, 5),
    28 => to_signed(1, 5),
    29 => to_signed(0, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(0, 5),
    33 => to_signed(-1, 5),
    34 => to_signed(-1, 5),
    35 => to_signed(-2, 5),
    36 => to_signed(-2, 5),
    37 => to_signed(-2, 5),
    38 => to_signed(-3, 5),
    39 => to_signed(-3, 5),
    40 => to_signed(-3, 5),
    41 => to_signed(-4, 5),
    42 => to_signed(-4, 5),
    43 => to_signed(-5, 5),
    44 => to_signed(-5, 5),
    45 => to_signed(-5, 5),
    46 => to_signed(-6, 5),
    47 => to_signed(-6, 5),
    48 => to_signed(-6, 5),
    49 => to_signed(-6, 5),
    50 => to_signed(-7, 5),
    51 => to_signed(-7, 5),
    52 => to_signed(-7, 5),
    53 => to_signed(-8, 5),
    54 => to_signed(-8, 5),
    55 => to_signed(-8, 5),
    56 => to_signed(-9, 5),
    57 => to_signed(-9, 5),
    58 => to_signed(-10, 5),
    59 => to_signed(-10, 5),
    60 => to_signed(-10, 5),
    61 => to_signed(-11, 5),
    62 => to_signed(-11, 5),
    63 => to_signed(-12, 5)
  );

  constant LUT_0_15_6_DATA : lut_array_t_0 := (
    0 => to_signed(-2, 5),
    1 => to_signed(-2, 5),
    2 => to_signed(-2, 5),
    3 => to_signed(-2, 5),
    4 => to_signed(-3, 5),
    5 => to_signed(-3, 5),
    6 => to_signed(-3, 5),
    7 => to_signed(-4, 5),
    8 => to_signed(-4, 5),
    9 => to_signed(-4, 5),
    10 => to_signed(-5, 5),
    11 => to_signed(-5, 5),
    12 => to_signed(-5, 5),
    13 => to_signed(-5, 5),
    14 => to_signed(-5, 5),
    15 => to_signed(-5, 5),
    16 => to_signed(-5, 5),
    17 => to_signed(-4, 5),
    18 => to_signed(-4, 5),
    19 => to_signed(-4, 5),
    20 => to_signed(-3, 5),
    21 => to_signed(-3, 5),
    22 => to_signed(-2, 5),
    23 => to_signed(-2, 5),
    24 => to_signed(-2, 5),
    25 => to_signed(-1, 5),
    26 => to_signed(-1, 5),
    27 => to_signed(0, 5),
    28 => to_signed(0, 5),
    29 => to_signed(1, 5),
    30 => to_signed(1, 5),
    31 => to_signed(1, 5),
    32 => to_signed(2, 5),
    33 => to_signed(2, 5),
    34 => to_signed(2, 5),
    35 => to_signed(3, 5),
    36 => to_signed(3, 5),
    37 => to_signed(3, 5),
    38 => to_signed(4, 5),
    39 => to_signed(4, 5),
    40 => to_signed(4, 5),
    41 => to_signed(5, 5),
    42 => to_signed(5, 5),
    43 => to_signed(5, 5),
    44 => to_signed(5, 5),
    45 => to_signed(6, 5),
    46 => to_signed(6, 5),
    47 => to_signed(6, 5),
    48 => to_signed(7, 5),
    49 => to_signed(7, 5),
    50 => to_signed(7, 5),
    51 => to_signed(8, 5),
    52 => to_signed(8, 5),
    53 => to_signed(8, 5),
    54 => to_signed(9, 5),
    55 => to_signed(9, 5),
    56 => to_signed(10, 5),
    57 => to_signed(10, 5),
    58 => to_signed(11, 5),
    59 => to_signed(11, 5),
    60 => to_signed(12, 5),
    61 => to_signed(12, 5),
    62 => to_signed(13, 5),
    63 => to_signed(14, 5)
  );

  constant LUT_0_15_7_DATA : lut_array_t_0 := (
    0 => to_signed(3, 5),
    1 => to_signed(3, 5),
    2 => to_signed(4, 5),
    3 => to_signed(5, 5),
    4 => to_signed(5, 5),
    5 => to_signed(6, 5),
    6 => to_signed(7, 5),
    7 => to_signed(7, 5),
    8 => to_signed(8, 5),
    9 => to_signed(8, 5),
    10 => to_signed(8, 5),
    11 => to_signed(8, 5),
    12 => to_signed(9, 5),
    13 => to_signed(9, 5),
    14 => to_signed(9, 5),
    15 => to_signed(9, 5),
    16 => to_signed(9, 5),
    17 => to_signed(8, 5),
    18 => to_signed(8, 5),
    19 => to_signed(8, 5),
    20 => to_signed(7, 5),
    21 => to_signed(7, 5),
    22 => to_signed(6, 5),
    23 => to_signed(5, 5),
    24 => to_signed(5, 5),
    25 => to_signed(4, 5),
    26 => to_signed(3, 5),
    27 => to_signed(3, 5),
    28 => to_signed(2, 5),
    29 => to_signed(1, 5),
    30 => to_signed(0, 5),
    31 => to_signed(0, 5),
    32 => to_signed(-1, 5),
    33 => to_signed(-2, 5),
    34 => to_signed(-2, 5),
    35 => to_signed(-3, 5),
    36 => to_signed(-4, 5),
    37 => to_signed(-4, 5),
    38 => to_signed(-5, 5),
    39 => to_signed(-5, 5),
    40 => to_signed(-6, 5),
    41 => to_signed(-7, 5),
    42 => to_signed(-8, 5),
    43 => to_signed(-8, 5),
    44 => to_signed(-9, 5),
    45 => to_signed(-9, 5),
    46 => to_signed(-10, 5),
    47 => to_signed(-11, 5),
    48 => to_signed(-11, 5),
    49 => to_signed(-12, 5),
    50 => to_signed(-12, 5),
    51 => to_signed(-13, 5),
    52 => to_signed(-13, 5),
    53 => to_signed(-13, 5),
    54 => to_signed(-14, 5),
    55 => to_signed(-14, 5),
    56 => to_signed(-14, 5),
    57 => to_signed(-15, 5),
    58 => to_signed(-15, 5),
    59 => to_signed(-15, 5),
    60 => to_signed(-15, 5),
    61 => to_signed(-16, 5),
    62 => to_signed(-16, 5),
    63 => to_signed(-16, 5)
  );

  -- Layer 1
  subtype lut_output_t_1 is signed(7 downto 0);
  type lut_array_t_1 is array (0 to 31) of lut_output_t_1;


  constant LUT_1_0_0_DATA : lut_array_t_1 := (
    0 => to_signed(-47, 8),
    1 => to_signed(-46, 8),
    2 => to_signed(-44, 8),
    3 => to_signed(-42, 8),
    4 => to_signed(-40, 8),
    5 => to_signed(-37, 8),
    6 => to_signed(-34, 8),
    7 => to_signed(-30, 8),
    8 => to_signed(-27, 8),
    9 => to_signed(-25, 8),
    10 => to_signed(-22, 8),
    11 => to_signed(-19, 8),
    12 => to_signed(-17, 8),
    13 => to_signed(-15, 8),
    14 => to_signed(-12, 8),
    15 => to_signed(-10, 8),
    16 => to_signed(-8, 8),
    17 => to_signed(-6, 8),
    18 => to_signed(-3, 8),
    19 => to_signed(-1, 8),
    20 => to_signed(2, 8),
    21 => to_signed(4, 8),
    22 => to_signed(7, 8),
    23 => to_signed(10, 8),
    24 => to_signed(13, 8),
    25 => to_signed(17, 8),
    26 => to_signed(21, 8),
    27 => to_signed(25, 8),
    28 => to_signed(30, 8),
    29 => to_signed(34, 8),
    30 => to_signed(38, 8),
    31 => to_signed(42, 8)
  );

  constant LUT_1_0_1_DATA : lut_array_t_1 := (
    0 => to_signed(-36, 8),
    1 => to_signed(-33, 8),
    2 => to_signed(-30, 8),
    3 => to_signed(-26, 8),
    4 => to_signed(-22, 8),
    5 => to_signed(-18, 8),
    6 => to_signed(-14, 8),
    7 => to_signed(-10, 8),
    8 => to_signed(-6, 8),
    9 => to_signed(-3, 8),
    10 => to_signed(0, 8),
    11 => to_signed(2, 8),
    12 => to_signed(4, 8),
    13 => to_signed(6, 8),
    14 => to_signed(8, 8),
    15 => to_signed(9, 8),
    16 => to_signed(9, 8),
    17 => to_signed(10, 8),
    18 => to_signed(10, 8),
    19 => to_signed(9, 8),
    20 => to_signed(9, 8),
    21 => to_signed(8, 8),
    22 => to_signed(7, 8),
    23 => to_signed(6, 8),
    24 => to_signed(4, 8),
    25 => to_signed(3, 8),
    26 => to_signed(2, 8),
    27 => to_signed(1, 8),
    28 => to_signed(0, 8),
    29 => to_signed(-1, 8),
    30 => to_signed(-3, 8),
    31 => to_signed(-3, 8)
  );

  constant LUT_1_0_2_DATA : lut_array_t_1 := (
    0 => to_signed(23, 8),
    1 => to_signed(22, 8),
    2 => to_signed(21, 8),
    3 => to_signed(19, 8),
    4 => to_signed(18, 8),
    5 => to_signed(16, 8),
    6 => to_signed(14, 8),
    7 => to_signed(12, 8),
    8 => to_signed(10, 8),
    9 => to_signed(8, 8),
    10 => to_signed(6, 8),
    11 => to_signed(4, 8),
    12 => to_signed(1, 8),
    13 => to_signed(-1, 8),
    14 => to_signed(-3, 8),
    15 => to_signed(-5, 8),
    16 => to_signed(-7, 8),
    17 => to_signed(-8, 8),
    18 => to_signed(-10, 8),
    19 => to_signed(-11, 8),
    20 => to_signed(-13, 8),
    21 => to_signed(-14, 8),
    22 => to_signed(-15, 8),
    23 => to_signed(-17, 8),
    24 => to_signed(-19, 8),
    25 => to_signed(-21, 8),
    26 => to_signed(-24, 8),
    27 => to_signed(-26, 8),
    28 => to_signed(-29, 8),
    29 => to_signed(-32, 8),
    30 => to_signed(-35, 8),
    31 => to_signed(-38, 8)
  );

  constant LUT_1_0_3_DATA : lut_array_t_1 := (
    0 => to_signed(3, 8),
    1 => to_signed(4, 8),
    2 => to_signed(5, 8),
    3 => to_signed(5, 8),
    4 => to_signed(6, 8),
    5 => to_signed(6, 8),
    6 => to_signed(7, 8),
    7 => to_signed(7, 8),
    8 => to_signed(7, 8),
    9 => to_signed(7, 8),
    10 => to_signed(7, 8),
    11 => to_signed(7, 8),
    12 => to_signed(7, 8),
    13 => to_signed(7, 8),
    14 => to_signed(6, 8),
    15 => to_signed(6, 8),
    16 => to_signed(6, 8),
    17 => to_signed(5, 8),
    18 => to_signed(5, 8),
    19 => to_signed(4, 8),
    20 => to_signed(4, 8),
    21 => to_signed(3, 8),
    22 => to_signed(2, 8),
    23 => to_signed(1, 8),
    24 => to_signed(0, 8),
    25 => to_signed(-2, 8),
    26 => to_signed(-3, 8),
    27 => to_signed(-5, 8),
    28 => to_signed(-7, 8),
    29 => to_signed(-9, 8),
    30 => to_signed(-11, 8),
    31 => to_signed(-13, 8)
  );

  constant LUT_1_0_4_DATA : lut_array_t_1 := (
    0 => to_signed(-4, 8),
    1 => to_signed(-5, 8),
    2 => to_signed(-5, 8),
    3 => to_signed(-5, 8),
    4 => to_signed(-5, 8),
    5 => to_signed(-5, 8),
    6 => to_signed(-5, 8),
    7 => to_signed(-5, 8),
    8 => to_signed(-4, 8),
    9 => to_signed(-4, 8),
    10 => to_signed(-4, 8),
    11 => to_signed(-3, 8),
    12 => to_signed(-3, 8),
    13 => to_signed(-2, 8),
    14 => to_signed(-1, 8),
    15 => to_signed(-1, 8),
    16 => to_signed(0, 8),
    17 => to_signed(0, 8),
    18 => to_signed(1, 8),
    19 => to_signed(1, 8),
    20 => to_signed(2, 8),
    21 => to_signed(2, 8),
    22 => to_signed(2, 8),
    23 => to_signed(2, 8),
    24 => to_signed(2, 8),
    25 => to_signed(2, 8),
    26 => to_signed(2, 8),
    27 => to_signed(2, 8),
    28 => to_signed(2, 8),
    29 => to_signed(2, 8),
    30 => to_signed(2, 8),
    31 => to_signed(2, 8)
  );

  constant LUT_1_1_0_DATA : lut_array_t_1 := (
    0 => to_signed(-10, 8),
    1 => to_signed(-10, 8),
    2 => to_signed(-10, 8),
    3 => to_signed(-10, 8),
    4 => to_signed(-11, 8),
    5 => to_signed(-11, 8),
    6 => to_signed(-11, 8),
    7 => to_signed(-10, 8),
    8 => to_signed(-10, 8),
    9 => to_signed(-10, 8),
    10 => to_signed(-9, 8),
    11 => to_signed(-9, 8),
    12 => to_signed(-8, 8),
    13 => to_signed(-7, 8),
    14 => to_signed(-6, 8),
    15 => to_signed(-5, 8),
    16 => to_signed(-4, 8),
    17 => to_signed(-3, 8),
    18 => to_signed(-2, 8),
    19 => to_signed(0, 8),
    20 => to_signed(1, 8),
    21 => to_signed(3, 8),
    22 => to_signed(4, 8),
    23 => to_signed(6, 8),
    24 => to_signed(8, 8),
    25 => to_signed(9, 8),
    26 => to_signed(11, 8),
    27 => to_signed(13, 8),
    28 => to_signed(14, 8),
    29 => to_signed(16, 8),
    30 => to_signed(17, 8),
    31 => to_signed(19, 8)
  );

  constant LUT_1_1_1_DATA : lut_array_t_1 := (
    0 => to_signed(4, 8),
    1 => to_signed(4, 8),
    2 => to_signed(3, 8),
    3 => to_signed(3, 8),
    4 => to_signed(3, 8),
    5 => to_signed(2, 8),
    6 => to_signed(2, 8),
    7 => to_signed(1, 8),
    8 => to_signed(1, 8),
    9 => to_signed(0, 8),
    10 => to_signed(-1, 8),
    11 => to_signed(-1, 8),
    12 => to_signed(-2, 8),
    13 => to_signed(-2, 8),
    14 => to_signed(-2, 8),
    15 => to_signed(-2, 8),
    16 => to_signed(-2, 8),
    17 => to_signed(-2, 8),
    18 => to_signed(-1, 8),
    19 => to_signed(-1, 8),
    20 => to_signed(0, 8),
    21 => to_signed(1, 8),
    22 => to_signed(1, 8),
    23 => to_signed(2, 8),
    24 => to_signed(3, 8),
    25 => to_signed(3, 8),
    26 => to_signed(3, 8),
    27 => to_signed(4, 8),
    28 => to_signed(4, 8),
    29 => to_signed(4, 8),
    30 => to_signed(4, 8),
    31 => to_signed(3, 8)
  );

  constant LUT_1_1_2_DATA : lut_array_t_1 := (
    0 => to_signed(-46, 8),
    1 => to_signed(-46, 8),
    2 => to_signed(-44, 8),
    3 => to_signed(-42, 8),
    4 => to_signed(-39, 8),
    5 => to_signed(-35, 8),
    6 => to_signed(-31, 8),
    7 => to_signed(-27, 8),
    8 => to_signed(-22, 8),
    9 => to_signed(-17, 8),
    10 => to_signed(-12, 8),
    11 => to_signed(-8, 8),
    12 => to_signed(-3, 8),
    13 => to_signed(1, 8),
    14 => to_signed(5, 8),
    15 => to_signed(8, 8),
    16 => to_signed(10, 8),
    17 => to_signed(11, 8),
    18 => to_signed(12, 8),
    19 => to_signed(12, 8),
    20 => to_signed(11, 8),
    21 => to_signed(9, 8),
    22 => to_signed(7, 8),
    23 => to_signed(5, 8),
    24 => to_signed(2, 8),
    25 => to_signed(-1, 8),
    26 => to_signed(-4, 8),
    27 => to_signed(-7, 8),
    28 => to_signed(-10, 8),
    29 => to_signed(-13, 8),
    30 => to_signed(-15, 8),
    31 => to_signed(-17, 8)
  );

  constant LUT_1_1_3_DATA : lut_array_t_1 := (
    0 => to_signed(-8, 8),
    1 => to_signed(-5, 8),
    2 => to_signed(-3, 8),
    3 => to_signed(0, 8),
    4 => to_signed(3, 8),
    5 => to_signed(5, 8),
    6 => to_signed(8, 8),
    7 => to_signed(9, 8),
    8 => to_signed(11, 8),
    9 => to_signed(11, 8),
    10 => to_signed(11, 8),
    11 => to_signed(11, 8),
    12 => to_signed(11, 8),
    13 => to_signed(10, 8),
    14 => to_signed(9, 8),
    15 => to_signed(8, 8),
    16 => to_signed(6, 8),
    17 => to_signed(5, 8),
    18 => to_signed(3, 8),
    19 => to_signed(2, 8),
    20 => to_signed(0, 8),
    21 => to_signed(-1, 8),
    22 => to_signed(-3, 8),
    23 => to_signed(-4, 8),
    24 => to_signed(-6, 8),
    25 => to_signed(-7, 8),
    26 => to_signed(-9, 8),
    27 => to_signed(-10, 8),
    28 => to_signed(-11, 8),
    29 => to_signed(-12, 8),
    30 => to_signed(-13, 8),
    31 => to_signed(-14, 8)
  );

  constant LUT_1_1_4_DATA : lut_array_t_1 := (
    0 => to_signed(17, 8),
    1 => to_signed(16, 8),
    2 => to_signed(16, 8),
    3 => to_signed(15, 8),
    4 => to_signed(14, 8),
    5 => to_signed(13, 8),
    6 => to_signed(12, 8),
    7 => to_signed(10, 8),
    8 => to_signed(9, 8),
    9 => to_signed(7, 8),
    10 => to_signed(5, 8),
    11 => to_signed(3, 8),
    12 => to_signed(1, 8),
    13 => to_signed(-2, 8),
    14 => to_signed(-4, 8),
    15 => to_signed(-6, 8),
    16 => to_signed(-8, 8),
    17 => to_signed(-9, 8),
    18 => to_signed(-11, 8),
    19 => to_signed(-13, 8),
    20 => to_signed(-14, 8),
    21 => to_signed(-15, 8),
    22 => to_signed(-16, 8),
    23 => to_signed(-17, 8),
    24 => to_signed(-18, 8),
    25 => to_signed(-18, 8),
    26 => to_signed(-18, 8),
    27 => to_signed(-19, 8),
    28 => to_signed(-19, 8),
    29 => to_signed(-18, 8),
    30 => to_signed(-18, 8),
    31 => to_signed(-18, 8)
  );

  constant LUT_1_2_0_DATA : lut_array_t_1 := (
    0 => to_signed(-28, 8),
    1 => to_signed(-27, 8),
    2 => to_signed(-26, 8),
    3 => to_signed(-25, 8),
    4 => to_signed(-25, 8),
    5 => to_signed(-24, 8),
    6 => to_signed(-23, 8),
    7 => to_signed(-22, 8),
    8 => to_signed(-22, 8),
    9 => to_signed(-21, 8),
    10 => to_signed(-21, 8),
    11 => to_signed(-20, 8),
    12 => to_signed(-19, 8),
    13 => to_signed(-18, 8),
    14 => to_signed(-17, 8),
    15 => to_signed(-16, 8),
    16 => to_signed(-14, 8),
    17 => to_signed(-11, 8),
    18 => to_signed(-8, 8),
    19 => to_signed(-5, 8),
    20 => to_signed(-1, 8),
    21 => to_signed(3, 8),
    22 => to_signed(8, 8),
    23 => to_signed(13, 8),
    24 => to_signed(18, 8),
    25 => to_signed(24, 8),
    26 => to_signed(31, 8),
    27 => to_signed(37, 8),
    28 => to_signed(44, 8),
    29 => to_signed(51, 8),
    30 => to_signed(57, 8),
    31 => to_signed(64, 8)
  );

  constant LUT_1_2_1_DATA : lut_array_t_1 := (
    0 => to_signed(27, 8),
    1 => to_signed(26, 8),
    2 => to_signed(25, 8),
    3 => to_signed(24, 8),
    4 => to_signed(23, 8),
    5 => to_signed(21, 8),
    6 => to_signed(19, 8),
    7 => to_signed(17, 8),
    8 => to_signed(15, 8),
    9 => to_signed(12, 8),
    10 => to_signed(10, 8),
    11 => to_signed(7, 8),
    12 => to_signed(4, 8),
    13 => to_signed(2, 8),
    14 => to_signed(-1, 8),
    15 => to_signed(-3, 8),
    16 => to_signed(-5, 8),
    17 => to_signed(-7, 8),
    18 => to_signed(-9, 8),
    19 => to_signed(-10, 8),
    20 => to_signed(-12, 8),
    21 => to_signed(-13, 8),
    22 => to_signed(-14, 8),
    23 => to_signed(-16, 8),
    24 => to_signed(-17, 8),
    25 => to_signed(-19, 8),
    26 => to_signed(-20, 8),
    27 => to_signed(-22, 8),
    28 => to_signed(-24, 8),
    29 => to_signed(-26, 8),
    30 => to_signed(-29, 8),
    31 => to_signed(-31, 8)
  );

  constant LUT_1_2_2_DATA : lut_array_t_1 := (
    0 => to_signed(-11, 8),
    1 => to_signed(-10, 8),
    2 => to_signed(-9, 8),
    3 => to_signed(-8, 8),
    4 => to_signed(-6, 8),
    5 => to_signed(-5, 8),
    6 => to_signed(-4, 8),
    7 => to_signed(-2, 8),
    8 => to_signed(-1, 8),
    9 => to_signed(1, 8),
    10 => to_signed(2, 8),
    11 => to_signed(4, 8),
    12 => to_signed(5, 8),
    13 => to_signed(6, 8),
    14 => to_signed(7, 8),
    15 => to_signed(7, 8),
    16 => to_signed(7, 8),
    17 => to_signed(7, 8),
    18 => to_signed(6, 8),
    19 => to_signed(4, 8),
    20 => to_signed(3, 8),
    21 => to_signed(1, 8),
    22 => to_signed(-2, 8),
    23 => to_signed(-5, 8),
    24 => to_signed(-8, 8),
    25 => to_signed(-12, 8),
    26 => to_signed(-16, 8),
    27 => to_signed(-20, 8),
    28 => to_signed(-24, 8),
    29 => to_signed(-29, 8),
    30 => to_signed(-32, 8),
    31 => to_signed(-36, 8)
  );

  constant LUT_1_2_3_DATA : lut_array_t_1 := (
    0 => to_signed(-7, 8),
    1 => to_signed(-7, 8),
    2 => to_signed(-6, 8),
    3 => to_signed(-5, 8),
    4 => to_signed(-4, 8),
    5 => to_signed(-3, 8),
    6 => to_signed(-2, 8),
    7 => to_signed(0, 8),
    8 => to_signed(1, 8),
    9 => to_signed(2, 8),
    10 => to_signed(3, 8),
    11 => to_signed(4, 8),
    12 => to_signed(6, 8),
    13 => to_signed(7, 8),
    14 => to_signed(8, 8),
    15 => to_signed(9, 8),
    16 => to_signed(10, 8),
    17 => to_signed(10, 8),
    18 => to_signed(11, 8),
    19 => to_signed(11, 8),
    20 => to_signed(10, 8),
    21 => to_signed(10, 8),
    22 => to_signed(8, 8),
    23 => to_signed(6, 8),
    24 => to_signed(3, 8),
    25 => to_signed(0, 8),
    26 => to_signed(-5, 8),
    27 => to_signed(-10, 8),
    28 => to_signed(-15, 8),
    29 => to_signed(-21, 8),
    30 => to_signed(-26, 8),
    31 => to_signed(-31, 8)
  );

  constant LUT_1_2_4_DATA : lut_array_t_1 := (
    0 => to_signed(5, 8),
    1 => to_signed(6, 8),
    2 => to_signed(7, 8),
    3 => to_signed(7, 8),
    4 => to_signed(8, 8),
    5 => to_signed(8, 8),
    6 => to_signed(8, 8),
    7 => to_signed(8, 8),
    8 => to_signed(8, 8),
    9 => to_signed(7, 8),
    10 => to_signed(7, 8),
    11 => to_signed(6, 8),
    12 => to_signed(5, 8),
    13 => to_signed(4, 8),
    14 => to_signed(3, 8),
    15 => to_signed(2, 8),
    16 => to_signed(1, 8),
    17 => to_signed(0, 8),
    18 => to_signed(-1, 8),
    19 => to_signed(-2, 8),
    20 => to_signed(-3, 8),
    21 => to_signed(-4, 8),
    22 => to_signed(-4, 8),
    23 => to_signed(-5, 8),
    24 => to_signed(-6, 8),
    25 => to_signed(-6, 8),
    26 => to_signed(-7, 8),
    27 => to_signed(-8, 8),
    28 => to_signed(-8, 8),
    29 => to_signed(-9, 8),
    30 => to_signed(-10, 8),
    31 => to_signed(-10, 8)
  );

  constant LUT_1_3_0_DATA : lut_array_t_1 := (
    0 => to_signed(-25, 8),
    1 => to_signed(-23, 8),
    2 => to_signed(-21, 8),
    3 => to_signed(-19, 8),
    4 => to_signed(-17, 8),
    5 => to_signed(-14, 8),
    6 => to_signed(-12, 8),
    7 => to_signed(-9, 8),
    8 => to_signed(-7, 8),
    9 => to_signed(-5, 8),
    10 => to_signed(-3, 8),
    11 => to_signed(-1, 8),
    12 => to_signed(1, 8),
    13 => to_signed(2, 8),
    14 => to_signed(3, 8),
    15 => to_signed(4, 8),
    16 => to_signed(5, 8),
    17 => to_signed(6, 8),
    18 => to_signed(6, 8),
    19 => to_signed(6, 8),
    20 => to_signed(6, 8),
    21 => to_signed(6, 8),
    22 => to_signed(6, 8),
    23 => to_signed(6, 8),
    24 => to_signed(6, 8),
    25 => to_signed(6, 8),
    26 => to_signed(6, 8),
    27 => to_signed(6, 8),
    28 => to_signed(6, 8),
    29 => to_signed(6, 8),
    30 => to_signed(7, 8),
    31 => to_signed(7, 8)
  );

  constant LUT_1_3_1_DATA : lut_array_t_1 := (
    0 => to_signed(17, 8),
    1 => to_signed(16, 8),
    2 => to_signed(15, 8),
    3 => to_signed(13, 8),
    4 => to_signed(12, 8),
    5 => to_signed(11, 8),
    6 => to_signed(9, 8),
    7 => to_signed(8, 8),
    8 => to_signed(6, 8),
    9 => to_signed(5, 8),
    10 => to_signed(4, 8),
    11 => to_signed(2, 8),
    12 => to_signed(1, 8),
    13 => to_signed(0, 8),
    14 => to_signed(-1, 8),
    15 => to_signed(-2, 8),
    16 => to_signed(-4, 8),
    17 => to_signed(-5, 8),
    18 => to_signed(-6, 8),
    19 => to_signed(-7, 8),
    20 => to_signed(-8, 8),
    21 => to_signed(-8, 8),
    22 => to_signed(-9, 8),
    23 => to_signed(-10, 8),
    24 => to_signed(-11, 8),
    25 => to_signed(-12, 8),
    26 => to_signed(-13, 8),
    27 => to_signed(-14, 8),
    28 => to_signed(-16, 8),
    29 => to_signed(-16, 8),
    30 => to_signed(-17, 8),
    31 => to_signed(-18, 8)
  );

  constant LUT_1_3_2_DATA : lut_array_t_1 := (
    0 => to_signed(-1, 8),
    1 => to_signed(0, 8),
    2 => to_signed(1, 8),
    3 => to_signed(2, 8),
    4 => to_signed(3, 8),
    5 => to_signed(4, 8),
    6 => to_signed(5, 8),
    7 => to_signed(6, 8),
    8 => to_signed(6, 8),
    9 => to_signed(7, 8),
    10 => to_signed(7, 8),
    11 => to_signed(7, 8),
    12 => to_signed(6, 8),
    13 => to_signed(6, 8),
    14 => to_signed(5, 8),
    15 => to_signed(4, 8),
    16 => to_signed(3, 8),
    17 => to_signed(2, 8),
    18 => to_signed(1, 8),
    19 => to_signed(-1, 8),
    20 => to_signed(-3, 8),
    21 => to_signed(-5, 8),
    22 => to_signed(-6, 8),
    23 => to_signed(-8, 8),
    24 => to_signed(-10, 8),
    25 => to_signed(-12, 8),
    26 => to_signed(-14, 8),
    27 => to_signed(-15, 8),
    28 => to_signed(-17, 8),
    29 => to_signed(-18, 8),
    30 => to_signed(-19, 8),
    31 => to_signed(-20, 8)
  );

  constant LUT_1_3_3_DATA : lut_array_t_1 := (
    0 => to_signed(18, 8),
    1 => to_signed(17, 8),
    2 => to_signed(17, 8),
    3 => to_signed(17, 8),
    4 => to_signed(17, 8),
    5 => to_signed(16, 8),
    6 => to_signed(16, 8),
    7 => to_signed(15, 8),
    8 => to_signed(14, 8),
    9 => to_signed(13, 8),
    10 => to_signed(12, 8),
    11 => to_signed(11, 8),
    12 => to_signed(10, 8),
    13 => to_signed(8, 8),
    14 => to_signed(6, 8),
    15 => to_signed(4, 8),
    16 => to_signed(2, 8),
    17 => to_signed(0, 8),
    18 => to_signed(-2, 8),
    19 => to_signed(-5, 8),
    20 => to_signed(-7, 8),
    21 => to_signed(-10, 8),
    22 => to_signed(-12, 8),
    23 => to_signed(-15, 8),
    24 => to_signed(-17, 8),
    25 => to_signed(-19, 8),
    26 => to_signed(-21, 8),
    27 => to_signed(-23, 8),
    28 => to_signed(-25, 8),
    29 => to_signed(-27, 8),
    30 => to_signed(-29, 8),
    31 => to_signed(-30, 8)
  );

  constant LUT_1_3_4_DATA : lut_array_t_1 := (
    0 => to_signed(-64, 8),
    1 => to_signed(-63, 8),
    2 => to_signed(-62, 8),
    3 => to_signed(-60, 8),
    4 => to_signed(-57, 8),
    5 => to_signed(-54, 8),
    6 => to_signed(-51, 8),
    7 => to_signed(-47, 8),
    8 => to_signed(-43, 8),
    9 => to_signed(-39, 8),
    10 => to_signed(-35, 8),
    11 => to_signed(-30, 8),
    12 => to_signed(-26, 8),
    13 => to_signed(-22, 8),
    14 => to_signed(-17, 8),
    15 => to_signed(-13, 8),
    16 => to_signed(-9, 8),
    17 => to_signed(-5, 8),
    18 => to_signed(0, 8),
    19 => to_signed(4, 8),
    20 => to_signed(8, 8),
    21 => to_signed(11, 8),
    22 => to_signed(15, 8),
    23 => to_signed(19, 8),
    24 => to_signed(22, 8),
    25 => to_signed(25, 8),
    26 => to_signed(28, 8),
    27 => to_signed(31, 8),
    28 => to_signed(33, 8),
    29 => to_signed(36, 8),
    30 => to_signed(38, 8),
    31 => to_signed(40, 8)
  );

  constant LUT_1_4_0_DATA : lut_array_t_1 := (
    0 => to_signed(-30, 8),
    1 => to_signed(-31, 8),
    2 => to_signed(-32, 8),
    3 => to_signed(-32, 8),
    4 => to_signed(-32, 8),
    5 => to_signed(-31, 8),
    6 => to_signed(-31, 8),
    7 => to_signed(-30, 8),
    8 => to_signed(-28, 8),
    9 => to_signed(-27, 8),
    10 => to_signed(-25, 8),
    11 => to_signed(-23, 8),
    12 => to_signed(-21, 8),
    13 => to_signed(-18, 8),
    14 => to_signed(-16, 8),
    15 => to_signed(-13, 8),
    16 => to_signed(-11, 8),
    17 => to_signed(-8, 8),
    18 => to_signed(-5, 8),
    19 => to_signed(-3, 8),
    20 => to_signed(0, 8),
    21 => to_signed(2, 8),
    22 => to_signed(5, 8),
    23 => to_signed(7, 8),
    24 => to_signed(9, 8),
    25 => to_signed(10, 8),
    26 => to_signed(12, 8),
    27 => to_signed(13, 8),
    28 => to_signed(14, 8),
    29 => to_signed(15, 8),
    30 => to_signed(16, 8),
    31 => to_signed(16, 8)
  );

  constant LUT_1_4_1_DATA : lut_array_t_1 := (
    0 => to_signed(-15, 8),
    1 => to_signed(-15, 8),
    2 => to_signed(-14, 8),
    3 => to_signed(-13, 8),
    4 => to_signed(-12, 8),
    5 => to_signed(-11, 8),
    6 => to_signed(-9, 8),
    7 => to_signed(-8, 8),
    8 => to_signed(-6, 8),
    9 => to_signed(-5, 8),
    10 => to_signed(-3, 8),
    11 => to_signed(-2, 8),
    12 => to_signed(-1, 8),
    13 => to_signed(0, 8),
    14 => to_signed(1, 8),
    15 => to_signed(2, 8),
    16 => to_signed(2, 8),
    17 => to_signed(2, 8),
    18 => to_signed(2, 8),
    19 => to_signed(1, 8),
    20 => to_signed(0, 8),
    21 => to_signed(0, 8),
    22 => to_signed(-1, 8),
    23 => to_signed(-2, 8),
    24 => to_signed(-3, 8),
    25 => to_signed(-4, 8),
    26 => to_signed(-5, 8),
    27 => to_signed(-5, 8),
    28 => to_signed(-6, 8),
    29 => to_signed(-7, 8),
    30 => to_signed(-7, 8),
    31 => to_signed(-8, 8)
  );

  constant LUT_1_4_2_DATA : lut_array_t_1 := (
    0 => to_signed(11, 8),
    1 => to_signed(11, 8),
    2 => to_signed(12, 8),
    3 => to_signed(13, 8),
    4 => to_signed(14, 8),
    5 => to_signed(14, 8),
    6 => to_signed(14, 8),
    7 => to_signed(14, 8),
    8 => to_signed(14, 8),
    9 => to_signed(13, 8),
    10 => to_signed(12, 8),
    11 => to_signed(11, 8),
    12 => to_signed(9, 8),
    13 => to_signed(7, 8),
    14 => to_signed(5, 8),
    15 => to_signed(3, 8),
    16 => to_signed(0, 8),
    17 => to_signed(-2, 8),
    18 => to_signed(-5, 8),
    19 => to_signed(-8, 8),
    20 => to_signed(-11, 8),
    21 => to_signed(-14, 8),
    22 => to_signed(-17, 8),
    23 => to_signed(-19, 8),
    24 => to_signed(-22, 8),
    25 => to_signed(-24, 8),
    26 => to_signed(-26, 8),
    27 => to_signed(-27, 8),
    28 => to_signed(-28, 8),
    29 => to_signed(-29, 8),
    30 => to_signed(-30, 8),
    31 => to_signed(-31, 8)
  );

  constant LUT_1_4_3_DATA : lut_array_t_1 := (
    0 => to_signed(35, 8),
    1 => to_signed(34, 8),
    2 => to_signed(33, 8),
    3 => to_signed(31, 8),
    4 => to_signed(30, 8),
    5 => to_signed(28, 8),
    6 => to_signed(25, 8),
    7 => to_signed(23, 8),
    8 => to_signed(20, 8),
    9 => to_signed(18, 8),
    10 => to_signed(15, 8),
    11 => to_signed(12, 8),
    12 => to_signed(9, 8),
    13 => to_signed(6, 8),
    14 => to_signed(3, 8),
    15 => to_signed(0, 8),
    16 => to_signed(-3, 8),
    17 => to_signed(-6, 8),
    18 => to_signed(-8, 8),
    19 => to_signed(-11, 8),
    20 => to_signed(-14, 8),
    21 => to_signed(-16, 8),
    22 => to_signed(-19, 8),
    23 => to_signed(-22, 8),
    24 => to_signed(-25, 8),
    25 => to_signed(-28, 8),
    26 => to_signed(-31, 8),
    27 => to_signed(-35, 8),
    28 => to_signed(-38, 8),
    29 => to_signed(-42, 8),
    30 => to_signed(-45, 8),
    31 => to_signed(-49, 8)
  );

  constant LUT_1_4_4_DATA : lut_array_t_1 := (
    0 => to_signed(-36, 8),
    1 => to_signed(-35, 8),
    2 => to_signed(-32, 8),
    3 => to_signed(-29, 8),
    4 => to_signed(-25, 8),
    5 => to_signed(-22, 8),
    6 => to_signed(-18, 8),
    7 => to_signed(-13, 8),
    8 => to_signed(-10, 8),
    9 => to_signed(-6, 8),
    10 => to_signed(-3, 8),
    11 => to_signed(0, 8),
    12 => to_signed(3, 8),
    13 => to_signed(5, 8),
    14 => to_signed(7, 8),
    15 => to_signed(8, 8),
    16 => to_signed(9, 8),
    17 => to_signed(10, 8),
    18 => to_signed(9, 8),
    19 => to_signed(9, 8),
    20 => to_signed(8, 8),
    21 => to_signed(7, 8),
    22 => to_signed(5, 8),
    23 => to_signed(3, 8),
    24 => to_signed(2, 8),
    25 => to_signed(0, 8),
    26 => to_signed(-2, 8),
    27 => to_signed(-4, 8),
    28 => to_signed(-5, 8),
    29 => to_signed(-7, 8),
    30 => to_signed(-9, 8),
    31 => to_signed(-11, 8)
  );

  constant LUT_1_5_0_DATA : lut_array_t_1 := (
    0 => to_signed(9, 8),
    1 => to_signed(9, 8),
    2 => to_signed(10, 8),
    3 => to_signed(11, 8),
    4 => to_signed(11, 8),
    5 => to_signed(12, 8),
    6 => to_signed(12, 8),
    7 => to_signed(12, 8),
    8 => to_signed(12, 8),
    9 => to_signed(12, 8),
    10 => to_signed(11, 8),
    11 => to_signed(10, 8),
    12 => to_signed(9, 8),
    13 => to_signed(8, 8),
    14 => to_signed(7, 8),
    15 => to_signed(5, 8),
    16 => to_signed(4, 8),
    17 => to_signed(2, 8),
    18 => to_signed(1, 8),
    19 => to_signed(-1, 8),
    20 => to_signed(-3, 8),
    21 => to_signed(-4, 8),
    22 => to_signed(-6, 8),
    23 => to_signed(-7, 8),
    24 => to_signed(-9, 8),
    25 => to_signed(-10, 8),
    26 => to_signed(-11, 8),
    27 => to_signed(-13, 8),
    28 => to_signed(-14, 8),
    29 => to_signed(-15, 8),
    30 => to_signed(-16, 8),
    31 => to_signed(-17, 8)
  );

  constant LUT_1_5_1_DATA : lut_array_t_1 := (
    0 => to_signed(15, 8),
    1 => to_signed(14, 8),
    2 => to_signed(13, 8),
    3 => to_signed(12, 8),
    4 => to_signed(10, 8),
    5 => to_signed(9, 8),
    6 => to_signed(8, 8),
    7 => to_signed(6, 8),
    8 => to_signed(5, 8),
    9 => to_signed(3, 8),
    10 => to_signed(2, 8),
    11 => to_signed(0, 8),
    12 => to_signed(-1, 8),
    13 => to_signed(-3, 8),
    14 => to_signed(-4, 8),
    15 => to_signed(-4, 8),
    16 => to_signed(-5, 8),
    17 => to_signed(-5, 8),
    18 => to_signed(-5, 8),
    19 => to_signed(-5, 8),
    20 => to_signed(-4, 8),
    21 => to_signed(-3, 8),
    22 => to_signed(-3, 8),
    23 => to_signed(-2, 8),
    24 => to_signed(-1, 8),
    25 => to_signed(0, 8),
    26 => to_signed(1, 8),
    27 => to_signed(2, 8),
    28 => to_signed(3, 8),
    29 => to_signed(4, 8),
    30 => to_signed(5, 8),
    31 => to_signed(6, 8)
  );

  constant LUT_1_5_2_DATA : lut_array_t_1 := (
    0 => to_signed(-63, 8),
    1 => to_signed(-63, 8),
    2 => to_signed(-62, 8),
    3 => to_signed(-60, 8),
    4 => to_signed(-58, 8),
    5 => to_signed(-55, 8),
    6 => to_signed(-51, 8),
    7 => to_signed(-47, 8),
    8 => to_signed(-42, 8),
    9 => to_signed(-36, 8),
    10 => to_signed(-31, 8),
    11 => to_signed(-24, 8),
    12 => to_signed(-18, 8),
    13 => to_signed(-12, 8),
    14 => to_signed(-6, 8),
    15 => to_signed(0, 8),
    16 => to_signed(6, 8),
    17 => to_signed(11, 8),
    18 => to_signed(16, 8),
    19 => to_signed(20, 8),
    20 => to_signed(24, 8),
    21 => to_signed(27, 8),
    22 => to_signed(29, 8),
    23 => to_signed(31, 8),
    24 => to_signed(31, 8),
    25 => to_signed(32, 8),
    26 => to_signed(31, 8),
    27 => to_signed(30, 8),
    28 => to_signed(28, 8),
    29 => to_signed(26, 8),
    30 => to_signed(25, 8),
    31 => to_signed(23, 8)
  );

  constant LUT_1_5_3_DATA : lut_array_t_1 := (
    0 => to_signed(-13, 8),
    1 => to_signed(-7, 8),
    2 => to_signed(-1, 8),
    3 => to_signed(5, 8),
    4 => to_signed(10, 8),
    5 => to_signed(15, 8),
    6 => to_signed(19, 8),
    7 => to_signed(22, 8),
    8 => to_signed(24, 8),
    9 => to_signed(25, 8),
    10 => to_signed(25, 8),
    11 => to_signed(24, 8),
    12 => to_signed(22, 8),
    13 => to_signed(20, 8),
    14 => to_signed(17, 8),
    15 => to_signed(14, 8),
    16 => to_signed(10, 8),
    17 => to_signed(6, 8),
    18 => to_signed(1, 8),
    19 => to_signed(-3, 8),
    20 => to_signed(-7, 8),
    21 => to_signed(-11, 8),
    22 => to_signed(-15, 8),
    23 => to_signed(-18, 8),
    24 => to_signed(-20, 8),
    25 => to_signed(-22, 8),
    26 => to_signed(-22, 8),
    27 => to_signed(-22, 8),
    28 => to_signed(-22, 8),
    29 => to_signed(-21, 8),
    30 => to_signed(-20, 8),
    31 => to_signed(-19, 8)
  );

  constant LUT_1_5_4_DATA : lut_array_t_1 := (
    0 => to_signed(5, 8),
    1 => to_signed(4, 8),
    2 => to_signed(3, 8),
    3 => to_signed(2, 8),
    4 => to_signed(1, 8),
    5 => to_signed(0, 8),
    6 => to_signed(-1, 8),
    7 => to_signed(-2, 8),
    8 => to_signed(-2, 8),
    9 => to_signed(-3, 8),
    10 => to_signed(-3, 8),
    11 => to_signed(-3, 8),
    12 => to_signed(-3, 8),
    13 => to_signed(-3, 8),
    14 => to_signed(-3, 8),
    15 => to_signed(-3, 8),
    16 => to_signed(-3, 8),
    17 => to_signed(-3, 8),
    18 => to_signed(-3, 8),
    19 => to_signed(-2, 8),
    20 => to_signed(-2, 8),
    21 => to_signed(-2, 8),
    22 => to_signed(-2, 8),
    23 => to_signed(-2, 8),
    24 => to_signed(-1, 8),
    25 => to_signed(-1, 8),
    26 => to_signed(-1, 8),
    27 => to_signed(-1, 8),
    28 => to_signed(-1, 8),
    29 => to_signed(-1, 8),
    30 => to_signed(-2, 8),
    31 => to_signed(-2, 8)
  );

  constant LUT_1_6_0_DATA : lut_array_t_1 := (
    0 => to_signed(8, 8),
    1 => to_signed(8, 8),
    2 => to_signed(9, 8),
    3 => to_signed(9, 8),
    4 => to_signed(9, 8),
    5 => to_signed(9, 8),
    6 => to_signed(9, 8),
    7 => to_signed(8, 8),
    8 => to_signed(7, 8),
    9 => to_signed(6, 8),
    10 => to_signed(4, 8),
    11 => to_signed(2, 8),
    12 => to_signed(0, 8),
    13 => to_signed(-2, 8),
    14 => to_signed(-4, 8),
    15 => to_signed(-6, 8),
    16 => to_signed(-8, 8),
    17 => to_signed(-10, 8),
    18 => to_signed(-11, 8),
    19 => to_signed(-12, 8),
    20 => to_signed(-14, 8),
    21 => to_signed(-14, 8),
    22 => to_signed(-15, 8),
    23 => to_signed(-15, 8),
    24 => to_signed(-15, 8),
    25 => to_signed(-15, 8),
    26 => to_signed(-14, 8),
    27 => to_signed(-14, 8),
    28 => to_signed(-13, 8),
    29 => to_signed(-12, 8),
    30 => to_signed(-11, 8),
    31 => to_signed(-10, 8)
  );

  constant LUT_1_6_1_DATA : lut_array_t_1 := (
    0 => to_signed(2, 8),
    1 => to_signed(1, 8),
    2 => to_signed(1, 8),
    3 => to_signed(0, 8),
    4 => to_signed(-1, 8),
    5 => to_signed(-2, 8),
    6 => to_signed(-3, 8),
    7 => to_signed(-4, 8),
    8 => to_signed(-5, 8),
    9 => to_signed(-7, 8),
    10 => to_signed(-8, 8),
    11 => to_signed(-10, 8),
    12 => to_signed(-11, 8),
    13 => to_signed(-12, 8),
    14 => to_signed(-12, 8),
    15 => to_signed(-12, 8),
    16 => to_signed(-11, 8),
    17 => to_signed(-10, 8),
    18 => to_signed(-8, 8),
    19 => to_signed(-6, 8),
    20 => to_signed(-3, 8),
    21 => to_signed(0, 8),
    22 => to_signed(3, 8),
    23 => to_signed(6, 8),
    24 => to_signed(9, 8),
    25 => to_signed(11, 8),
    26 => to_signed(14, 8),
    27 => to_signed(16, 8),
    28 => to_signed(18, 8),
    29 => to_signed(19, 8),
    30 => to_signed(21, 8),
    31 => to_signed(22, 8)
  );

  constant LUT_1_6_2_DATA : lut_array_t_1 := (
    0 => to_signed(-6, 8),
    1 => to_signed(-6, 8),
    2 => to_signed(-6, 8),
    3 => to_signed(-6, 8),
    4 => to_signed(-5, 8),
    5 => to_signed(-4, 8),
    6 => to_signed(-3, 8),
    7 => to_signed(-2, 8),
    8 => to_signed(0, 8),
    9 => to_signed(2, 8),
    10 => to_signed(4, 8),
    11 => to_signed(6, 8),
    12 => to_signed(8, 8),
    13 => to_signed(9, 8),
    14 => to_signed(10, 8),
    15 => to_signed(10, 8),
    16 => to_signed(9, 8),
    17 => to_signed(8, 8),
    18 => to_signed(5, 8),
    19 => to_signed(2, 8),
    20 => to_signed(-2, 8),
    21 => to_signed(-7, 8),
    22 => to_signed(-12, 8),
    23 => to_signed(-17, 8),
    24 => to_signed(-23, 8),
    25 => to_signed(-28, 8),
    26 => to_signed(-34, 8),
    27 => to_signed(-39, 8),
    28 => to_signed(-44, 8),
    29 => to_signed(-48, 8),
    30 => to_signed(-52, 8),
    31 => to_signed(-56, 8)
  );

  constant LUT_1_6_3_DATA : lut_array_t_1 := (
    0 => to_signed(3, 8),
    1 => to_signed(3, 8),
    2 => to_signed(3, 8),
    3 => to_signed(3, 8),
    4 => to_signed(3, 8),
    5 => to_signed(3, 8),
    6 => to_signed(3, 8),
    7 => to_signed(4, 8),
    8 => to_signed(4, 8),
    9 => to_signed(5, 8),
    10 => to_signed(6, 8),
    11 => to_signed(7, 8),
    12 => to_signed(8, 8),
    13 => to_signed(9, 8),
    14 => to_signed(10, 8),
    15 => to_signed(11, 8),
    16 => to_signed(12, 8),
    17 => to_signed(12, 8),
    18 => to_signed(13, 8),
    19 => to_signed(12, 8),
    20 => to_signed(12, 8),
    21 => to_signed(10, 8),
    22 => to_signed(8, 8),
    23 => to_signed(5, 8),
    24 => to_signed(0, 8),
    25 => to_signed(-6, 8),
    26 => to_signed(-12, 8),
    27 => to_signed(-20, 8),
    28 => to_signed(-29, 8),
    29 => to_signed(-37, 8),
    30 => to_signed(-46, 8),
    31 => to_signed(-55, 8)
  );

  constant LUT_1_6_4_DATA : lut_array_t_1 := (
    0 => to_signed(-33, 8),
    1 => to_signed(-33, 8),
    2 => to_signed(-33, 8),
    3 => to_signed(-33, 8),
    4 => to_signed(-33, 8),
    5 => to_signed(-33, 8),
    6 => to_signed(-33, 8),
    7 => to_signed(-33, 8),
    8 => to_signed(-33, 8),
    9 => to_signed(-33, 8),
    10 => to_signed(-33, 8),
    11 => to_signed(-33, 8),
    12 => to_signed(-33, 8),
    13 => to_signed(-32, 8),
    14 => to_signed(-31, 8),
    15 => to_signed(-29, 8),
    16 => to_signed(-26, 8),
    17 => to_signed(-23, 8),
    18 => to_signed(-19, 8),
    19 => to_signed(-14, 8),
    20 => to_signed(-8, 8),
    21 => to_signed(-2, 8),
    22 => to_signed(3, 8),
    23 => to_signed(9, 8),
    24 => to_signed(15, 8),
    25 => to_signed(21, 8),
    26 => to_signed(26, 8),
    27 => to_signed(31, 8),
    28 => to_signed(36, 8),
    29 => to_signed(40, 8),
    30 => to_signed(44, 8),
    31 => to_signed(48, 8)
  );

  constant LUT_1_7_0_DATA : lut_array_t_1 := (
    0 => to_signed(10, 8),
    1 => to_signed(11, 8),
    2 => to_signed(12, 8),
    3 => to_signed(13, 8),
    4 => to_signed(14, 8),
    5 => to_signed(15, 8),
    6 => to_signed(16, 8),
    7 => to_signed(16, 8),
    8 => to_signed(16, 8),
    9 => to_signed(15, 8),
    10 => to_signed(15, 8),
    11 => to_signed(14, 8),
    12 => to_signed(12, 8),
    13 => to_signed(10, 8),
    14 => to_signed(8, 8),
    15 => to_signed(6, 8),
    16 => to_signed(4, 8),
    17 => to_signed(1, 8),
    18 => to_signed(-2, 8),
    19 => to_signed(-6, 8),
    20 => to_signed(-9, 8),
    21 => to_signed(-13, 8),
    22 => to_signed(-17, 8),
    23 => to_signed(-21, 8),
    24 => to_signed(-25, 8),
    25 => to_signed(-30, 8),
    26 => to_signed(-34, 8),
    27 => to_signed(-38, 8),
    28 => to_signed(-42, 8),
    29 => to_signed(-46, 8),
    30 => to_signed(-50, 8),
    31 => to_signed(-54, 8)
  );

  constant LUT_1_7_1_DATA : lut_array_t_1 := (
    0 => to_signed(14, 8),
    1 => to_signed(14, 8),
    2 => to_signed(14, 8),
    3 => to_signed(15, 8),
    4 => to_signed(15, 8),
    5 => to_signed(16, 8),
    6 => to_signed(16, 8),
    7 => to_signed(16, 8),
    8 => to_signed(16, 8),
    9 => to_signed(16, 8),
    10 => to_signed(16, 8),
    11 => to_signed(15, 8),
    12 => to_signed(15, 8),
    13 => to_signed(13, 8),
    14 => to_signed(12, 8),
    15 => to_signed(10, 8),
    16 => to_signed(8, 8),
    17 => to_signed(4, 8),
    18 => to_signed(1, 8),
    19 => to_signed(-3, 8),
    20 => to_signed(-8, 8),
    21 => to_signed(-12, 8),
    22 => to_signed(-18, 8),
    23 => to_signed(-23, 8),
    24 => to_signed(-28, 8),
    25 => to_signed(-34, 8),
    26 => to_signed(-40, 8),
    27 => to_signed(-46, 8),
    28 => to_signed(-52, 8),
    29 => to_signed(-57, 8),
    30 => to_signed(-63, 8),
    31 => to_signed(-68, 8)
  );

  constant LUT_1_7_2_DATA : lut_array_t_1 := (
    0 => to_signed(-28, 8),
    1 => to_signed(-27, 8),
    2 => to_signed(-27, 8),
    3 => to_signed(-26, 8),
    4 => to_signed(-25, 8),
    5 => to_signed(-24, 8),
    6 => to_signed(-22, 8),
    7 => to_signed(-21, 8),
    8 => to_signed(-19, 8),
    9 => to_signed(-17, 8),
    10 => to_signed(-15, 8),
    11 => to_signed(-13, 8),
    12 => to_signed(-11, 8),
    13 => to_signed(-9, 8),
    14 => to_signed(-7, 8),
    15 => to_signed(-5, 8),
    16 => to_signed(-2, 8),
    17 => to_signed(0, 8),
    18 => to_signed(3, 8),
    19 => to_signed(5, 8),
    20 => to_signed(7, 8),
    21 => to_signed(10, 8),
    22 => to_signed(12, 8),
    23 => to_signed(14, 8),
    24 => to_signed(16, 8),
    25 => to_signed(18, 8),
    26 => to_signed(20, 8),
    27 => to_signed(21, 8),
    28 => to_signed(23, 8),
    29 => to_signed(24, 8),
    30 => to_signed(25, 8),
    31 => to_signed(27, 8)
  );

  constant LUT_1_7_3_DATA : lut_array_t_1 := (
    0 => to_signed(-1, 8),
    1 => to_signed(-1, 8),
    2 => to_signed(-1, 8),
    3 => to_signed(-1, 8),
    4 => to_signed(-1, 8),
    5 => to_signed(0, 8),
    6 => to_signed(0, 8),
    7 => to_signed(0, 8),
    8 => to_signed(0, 8),
    9 => to_signed(0, 8),
    10 => to_signed(0, 8),
    11 => to_signed(0, 8),
    12 => to_signed(0, 8),
    13 => to_signed(0, 8),
    14 => to_signed(0, 8),
    15 => to_signed(0, 8),
    16 => to_signed(0, 8),
    17 => to_signed(0, 8),
    18 => to_signed(1, 8),
    19 => to_signed(1, 8),
    20 => to_signed(2, 8),
    21 => to_signed(3, 8),
    22 => to_signed(3, 8),
    23 => to_signed(4, 8),
    24 => to_signed(5, 8),
    25 => to_signed(6, 8),
    26 => to_signed(7, 8),
    27 => to_signed(8, 8),
    28 => to_signed(9, 8),
    29 => to_signed(10, 8),
    30 => to_signed(11, 8),
    31 => to_signed(11, 8)
  );

  constant LUT_1_7_4_DATA : lut_array_t_1 := (
    0 => to_signed(-27, 8),
    1 => to_signed(-28, 8),
    2 => to_signed(-28, 8),
    3 => to_signed(-29, 8),
    4 => to_signed(-28, 8),
    5 => to_signed(-28, 8),
    6 => to_signed(-27, 8),
    7 => to_signed(-26, 8),
    8 => to_signed(-24, 8),
    9 => to_signed(-22, 8),
    10 => to_signed(-20, 8),
    11 => to_signed(-17, 8),
    12 => to_signed(-15, 8),
    13 => to_signed(-12, 8),
    14 => to_signed(-9, 8),
    15 => to_signed(-6, 8),
    16 => to_signed(-3, 8),
    17 => to_signed(-1, 8),
    18 => to_signed(1, 8),
    19 => to_signed(3, 8),
    20 => to_signed(5, 8),
    21 => to_signed(6, 8),
    22 => to_signed(8, 8),
    23 => to_signed(9, 8),
    24 => to_signed(10, 8),
    25 => to_signed(11, 8),
    26 => to_signed(12, 8),
    27 => to_signed(13, 8),
    28 => to_signed(14, 8),
    29 => to_signed(15, 8),
    30 => to_signed(15, 8),
    31 => to_signed(16, 8)
  );
end package;