library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package PkgKAN is
  -- Model parameters
  constant N_INPUT  : positive := 128;
  constant N_OUTPUT : positive := 128;

  -- bitwidths
  constant INPUT_WIDTH : positive := 6;
  constant OUTPUT_WIDTH : positive := 6;

  subtype input_t  is unsigned(INPUT_WIDTH-1 downto 0);
  subtype output_t is signed(OUTPUT_WIDTH-1 downto 0);

  type input_vec_t  is array (0 to N_INPUT-1)  of input_t;
  type output_vec_t is array (0 to N_OUTPUT-1) of output_t;

  -- For summation
  constant SUM_WIDTH_0_0: positive := 6;
  subtype sum_t_0_0 is signed(SUM_WIDTH_0_0-1 downto 0);
  constant SUM_WIDTH_0_1: positive := 12;
  subtype sum_t_0_1 is signed(SUM_WIDTH_0_1-1 downto 0);
  constant SUM_WIDTH_0_2: positive := 6;
  subtype sum_t_0_2 is signed(SUM_WIDTH_0_2-1 downto 0);
  constant SUM_WIDTH_0_3: positive := 6;
  subtype sum_t_0_3 is signed(SUM_WIDTH_0_3-1 downto 0);
  constant SUM_WIDTH_0_4: positive := 13;
  subtype sum_t_0_4 is signed(SUM_WIDTH_0_4-1 downto 0);
  constant SUM_WIDTH_0_5: positive := 13;
  subtype sum_t_0_5 is signed(SUM_WIDTH_0_5-1 downto 0);
  constant SUM_WIDTH_0_6: positive := 6;
  subtype sum_t_0_6 is signed(SUM_WIDTH_0_6-1 downto 0);
  constant SUM_WIDTH_0_7: positive := 6;
  subtype sum_t_0_7 is signed(SUM_WIDTH_0_7-1 downto 0);
  constant SUM_WIDTH_1_0: positive := 6;
  subtype sum_t_1_0 is signed(SUM_WIDTH_1_0-1 downto 0);
  constant SUM_WIDTH_1_1: positive := 7;
  subtype sum_t_1_1 is signed(SUM_WIDTH_1_1-1 downto 0);
  constant SUM_WIDTH_1_2: positive := 6;
  subtype sum_t_1_2 is signed(SUM_WIDTH_1_2-1 downto 0);
  constant SUM_WIDTH_1_3: positive := 6;
  subtype sum_t_1_3 is signed(SUM_WIDTH_1_3-1 downto 0);
  constant SUM_WIDTH_1_4: positive := 7;
  subtype sum_t_1_4 is signed(SUM_WIDTH_1_4-1 downto 0);
  constant SUM_WIDTH_1_5: positive := 6;
  subtype sum_t_1_5 is signed(SUM_WIDTH_1_5-1 downto 0);
  constant SUM_WIDTH_1_6: positive := 7;
  subtype sum_t_1_6 is signed(SUM_WIDTH_1_6-1 downto 0);
  constant SUM_WIDTH_1_7: positive := 6;
  subtype sum_t_1_7 is signed(SUM_WIDTH_1_7-1 downto 0);
  constant SUM_WIDTH_2_0: positive := 7;
  subtype sum_t_2_0 is signed(SUM_WIDTH_2_0-1 downto 0);
  constant SUM_WIDTH_2_1: positive := 8;
  subtype sum_t_2_1 is signed(SUM_WIDTH_2_1-1 downto 0);
  constant SUM_WIDTH_2_2: positive := 6;
  subtype sum_t_2_2 is signed(SUM_WIDTH_2_2-1 downto 0);
  constant SUM_WIDTH_2_3: positive := 6;
  subtype sum_t_2_3 is signed(SUM_WIDTH_2_3-1 downto 0);
  constant SUM_WIDTH_2_4: positive := 8;
  subtype sum_t_2_4 is signed(SUM_WIDTH_2_4-1 downto 0);
  constant SUM_WIDTH_2_5: positive := 9;
  subtype sum_t_2_5 is signed(SUM_WIDTH_2_5-1 downto 0);
  constant SUM_WIDTH_2_6: positive := 9;
  subtype sum_t_2_6 is signed(SUM_WIDTH_2_6-1 downto 0);
  constant SUM_WIDTH_2_7: positive := 7;
  subtype sum_t_2_7 is signed(SUM_WIDTH_2_7-1 downto 0);
  constant SUM_WIDTH_3_0: positive := 9;
  subtype sum_t_3_0 is signed(SUM_WIDTH_3_0-1 downto 0);
  constant SUM_WIDTH_3_1: positive := 8;
  subtype sum_t_3_1 is signed(SUM_WIDTH_3_1-1 downto 0);
  constant SUM_WIDTH_3_2: positive := 7;
  subtype sum_t_3_2 is signed(SUM_WIDTH_3_2-1 downto 0);
  constant SUM_WIDTH_3_3: positive := 9;
  subtype sum_t_3_3 is signed(SUM_WIDTH_3_3-1 downto 0);
  constant SUM_WIDTH_3_4: positive := 8;
  subtype sum_t_3_4 is signed(SUM_WIDTH_3_4-1 downto 0);
  constant SUM_WIDTH_3_5: positive := 9;
  subtype sum_t_3_5 is signed(SUM_WIDTH_3_5-1 downto 0);
  constant SUM_WIDTH_3_6: positive := 8;
  subtype sum_t_3_6 is signed(SUM_WIDTH_3_6-1 downto 0);
  constant SUM_WIDTH_3_7: positive := 9;
  subtype sum_t_3_7 is signed(SUM_WIDTH_3_7-1 downto 0);
  constant SUM_WIDTH_3_8: positive := 9;
  subtype sum_t_3_8 is signed(SUM_WIDTH_3_8-1 downto 0);
  constant SUM_WIDTH_3_9: positive := 9;
  subtype sum_t_3_9 is signed(SUM_WIDTH_3_9-1 downto 0);
  constant SUM_WIDTH_3_10: positive := 8;
  subtype sum_t_3_10 is signed(SUM_WIDTH_3_10-1 downto 0);
  constant SUM_WIDTH_3_11: positive := 9;
  subtype sum_t_3_11 is signed(SUM_WIDTH_3_11-1 downto 0);
  constant SUM_WIDTH_3_12: positive := 9;
  subtype sum_t_3_12 is signed(SUM_WIDTH_3_12-1 downto 0);
  constant SUM_WIDTH_3_13: positive := 9;
  subtype sum_t_3_13 is signed(SUM_WIDTH_3_13-1 downto 0);
  constant SUM_WIDTH_3_14: positive := 8;
  subtype sum_t_3_14 is signed(SUM_WIDTH_3_14-1 downto 0);
  constant SUM_WIDTH_3_15: positive := 8;
  subtype sum_t_3_15 is signed(SUM_WIDTH_3_15-1 downto 0);
  constant SUM_WIDTH_3_16: positive := 9;
  subtype sum_t_3_16 is signed(SUM_WIDTH_3_16-1 downto 0);
  constant SUM_WIDTH_3_17: positive := 8;
  subtype sum_t_3_17 is signed(SUM_WIDTH_3_17-1 downto 0);
  constant SUM_WIDTH_3_18: positive := 8;
  subtype sum_t_3_18 is signed(SUM_WIDTH_3_18-1 downto 0);
  constant SUM_WIDTH_3_19: positive := 8;
  subtype sum_t_3_19 is signed(SUM_WIDTH_3_19-1 downto 0);
  constant SUM_WIDTH_3_20: positive := 9;
  subtype sum_t_3_20 is signed(SUM_WIDTH_3_20-1 downto 0);
  constant SUM_WIDTH_3_21: positive := 8;
  subtype sum_t_3_21 is signed(SUM_WIDTH_3_21-1 downto 0);
  constant SUM_WIDTH_3_22: positive := 7;
  subtype sum_t_3_22 is signed(SUM_WIDTH_3_22-1 downto 0);
  constant SUM_WIDTH_3_23: positive := 8;
  subtype sum_t_3_23 is signed(SUM_WIDTH_3_23-1 downto 0);
  constant SUM_WIDTH_3_24: positive := 9;
  subtype sum_t_3_24 is signed(SUM_WIDTH_3_24-1 downto 0);
  constant SUM_WIDTH_3_25: positive := 9;
  subtype sum_t_3_25 is signed(SUM_WIDTH_3_25-1 downto 0);
  constant SUM_WIDTH_3_26: positive := 8;
  subtype sum_t_3_26 is signed(SUM_WIDTH_3_26-1 downto 0);
  constant SUM_WIDTH_3_27: positive := 9;
  subtype sum_t_3_27 is signed(SUM_WIDTH_3_27-1 downto 0);
  constant SUM_WIDTH_3_28: positive := 9;
  subtype sum_t_3_28 is signed(SUM_WIDTH_3_28-1 downto 0);
  constant SUM_WIDTH_3_29: positive := 9;
  subtype sum_t_3_29 is signed(SUM_WIDTH_3_29-1 downto 0);
  constant SUM_WIDTH_3_30: positive := 9;
  subtype sum_t_3_30 is signed(SUM_WIDTH_3_30-1 downto 0);
  constant SUM_WIDTH_3_31: positive := 9;
  subtype sum_t_3_31 is signed(SUM_WIDTH_3_31-1 downto 0);
  constant SUM_WIDTH_3_32: positive := 9;
  subtype sum_t_3_32 is signed(SUM_WIDTH_3_32-1 downto 0);
  constant SUM_WIDTH_3_33: positive := 9;
  subtype sum_t_3_33 is signed(SUM_WIDTH_3_33-1 downto 0);
  constant SUM_WIDTH_3_34: positive := 9;
  subtype sum_t_3_34 is signed(SUM_WIDTH_3_34-1 downto 0);
  constant SUM_WIDTH_3_35: positive := 9;
  subtype sum_t_3_35 is signed(SUM_WIDTH_3_35-1 downto 0);
  constant SUM_WIDTH_3_36: positive := 9;
  subtype sum_t_3_36 is signed(SUM_WIDTH_3_36-1 downto 0);
  constant SUM_WIDTH_3_37: positive := 9;
  subtype sum_t_3_37 is signed(SUM_WIDTH_3_37-1 downto 0);
  constant SUM_WIDTH_3_38: positive := 8;
  subtype sum_t_3_38 is signed(SUM_WIDTH_3_38-1 downto 0);
  constant SUM_WIDTH_3_39: positive := 9;
  subtype sum_t_3_39 is signed(SUM_WIDTH_3_39-1 downto 0);
  constant SUM_WIDTH_3_40: positive := 9;
  subtype sum_t_3_40 is signed(SUM_WIDTH_3_40-1 downto 0);
  constant SUM_WIDTH_3_41: positive := 9;
  subtype sum_t_3_41 is signed(SUM_WIDTH_3_41-1 downto 0);
  constant SUM_WIDTH_3_42: positive := 9;
  subtype sum_t_3_42 is signed(SUM_WIDTH_3_42-1 downto 0);
  constant SUM_WIDTH_3_43: positive := 9;
  subtype sum_t_3_43 is signed(SUM_WIDTH_3_43-1 downto 0);
  constant SUM_WIDTH_3_44: positive := 9;
  subtype sum_t_3_44 is signed(SUM_WIDTH_3_44-1 downto 0);
  constant SUM_WIDTH_3_45: positive := 8;
  subtype sum_t_3_45 is signed(SUM_WIDTH_3_45-1 downto 0);
  constant SUM_WIDTH_3_46: positive := 9;
  subtype sum_t_3_46 is signed(SUM_WIDTH_3_46-1 downto 0);
  constant SUM_WIDTH_3_47: positive := 9;
  subtype sum_t_3_47 is signed(SUM_WIDTH_3_47-1 downto 0);
  constant SUM_WIDTH_3_48: positive := 9;
  subtype sum_t_3_48 is signed(SUM_WIDTH_3_48-1 downto 0);
  constant SUM_WIDTH_3_49: positive := 8;
  subtype sum_t_3_49 is signed(SUM_WIDTH_3_49-1 downto 0);
  constant SUM_WIDTH_3_50: positive := 9;
  subtype sum_t_3_50 is signed(SUM_WIDTH_3_50-1 downto 0);
  constant SUM_WIDTH_3_51: positive := 9;
  subtype sum_t_3_51 is signed(SUM_WIDTH_3_51-1 downto 0);
  constant SUM_WIDTH_3_52: positive := 9;
  subtype sum_t_3_52 is signed(SUM_WIDTH_3_52-1 downto 0);
  constant SUM_WIDTH_3_53: positive := 9;
  subtype sum_t_3_53 is signed(SUM_WIDTH_3_53-1 downto 0);
  constant SUM_WIDTH_3_54: positive := 8;
  subtype sum_t_3_54 is signed(SUM_WIDTH_3_54-1 downto 0);
  constant SUM_WIDTH_3_55: positive := 9;
  subtype sum_t_3_55 is signed(SUM_WIDTH_3_55-1 downto 0);
  constant SUM_WIDTH_3_56: positive := 9;
  subtype sum_t_3_56 is signed(SUM_WIDTH_3_56-1 downto 0);
  constant SUM_WIDTH_3_57: positive := 8;
  subtype sum_t_3_57 is signed(SUM_WIDTH_3_57-1 downto 0);
  constant SUM_WIDTH_3_58: positive := 9;
  subtype sum_t_3_58 is signed(SUM_WIDTH_3_58-1 downto 0);
  constant SUM_WIDTH_3_59: positive := 8;
  subtype sum_t_3_59 is signed(SUM_WIDTH_3_59-1 downto 0);
  constant SUM_WIDTH_3_60: positive := 9;
  subtype sum_t_3_60 is signed(SUM_WIDTH_3_60-1 downto 0);
  constant SUM_WIDTH_3_61: positive := 9;
  subtype sum_t_3_61 is signed(SUM_WIDTH_3_61-1 downto 0);
  constant SUM_WIDTH_3_62: positive := 8;
  subtype sum_t_3_62 is signed(SUM_WIDTH_3_62-1 downto 0);
  constant SUM_WIDTH_3_63: positive := 8;
  subtype sum_t_3_63 is signed(SUM_WIDTH_3_63-1 downto 0);
  constant SUM_WIDTH_3_64: positive := 9;
  subtype sum_t_3_64 is signed(SUM_WIDTH_3_64-1 downto 0);
  constant SUM_WIDTH_3_65: positive := 8;
  subtype sum_t_3_65 is signed(SUM_WIDTH_3_65-1 downto 0);
  constant SUM_WIDTH_3_66: positive := 9;
  subtype sum_t_3_66 is signed(SUM_WIDTH_3_66-1 downto 0);
  constant SUM_WIDTH_3_67: positive := 8;
  subtype sum_t_3_67 is signed(SUM_WIDTH_3_67-1 downto 0);
  constant SUM_WIDTH_3_68: positive := 9;
  subtype sum_t_3_68 is signed(SUM_WIDTH_3_68-1 downto 0);
  constant SUM_WIDTH_3_69: positive := 9;
  subtype sum_t_3_69 is signed(SUM_WIDTH_3_69-1 downto 0);
  constant SUM_WIDTH_3_70: positive := 9;
  subtype sum_t_3_70 is signed(SUM_WIDTH_3_70-1 downto 0);
  constant SUM_WIDTH_3_71: positive := 9;
  subtype sum_t_3_71 is signed(SUM_WIDTH_3_71-1 downto 0);
  constant SUM_WIDTH_3_72: positive := 9;
  subtype sum_t_3_72 is signed(SUM_WIDTH_3_72-1 downto 0);
  constant SUM_WIDTH_3_73: positive := 8;
  subtype sum_t_3_73 is signed(SUM_WIDTH_3_73-1 downto 0);
  constant SUM_WIDTH_3_74: positive := 9;
  subtype sum_t_3_74 is signed(SUM_WIDTH_3_74-1 downto 0);
  constant SUM_WIDTH_3_75: positive := 8;
  subtype sum_t_3_75 is signed(SUM_WIDTH_3_75-1 downto 0);
  constant SUM_WIDTH_3_76: positive := 9;
  subtype sum_t_3_76 is signed(SUM_WIDTH_3_76-1 downto 0);
  constant SUM_WIDTH_3_77: positive := 9;
  subtype sum_t_3_77 is signed(SUM_WIDTH_3_77-1 downto 0);
  constant SUM_WIDTH_3_78: positive := 9;
  subtype sum_t_3_78 is signed(SUM_WIDTH_3_78-1 downto 0);
  constant SUM_WIDTH_3_79: positive := 9;
  subtype sum_t_3_79 is signed(SUM_WIDTH_3_79-1 downto 0);
  constant SUM_WIDTH_3_80: positive := 9;
  subtype sum_t_3_80 is signed(SUM_WIDTH_3_80-1 downto 0);
  constant SUM_WIDTH_3_81: positive := 8;
  subtype sum_t_3_81 is signed(SUM_WIDTH_3_81-1 downto 0);
  constant SUM_WIDTH_3_82: positive := 9;
  subtype sum_t_3_82 is signed(SUM_WIDTH_3_82-1 downto 0);
  constant SUM_WIDTH_3_83: positive := 9;
  subtype sum_t_3_83 is signed(SUM_WIDTH_3_83-1 downto 0);
  constant SUM_WIDTH_3_84: positive := 8;
  subtype sum_t_3_84 is signed(SUM_WIDTH_3_84-1 downto 0);
  constant SUM_WIDTH_3_85: positive := 9;
  subtype sum_t_3_85 is signed(SUM_WIDTH_3_85-1 downto 0);
  constant SUM_WIDTH_3_86: positive := 9;
  subtype sum_t_3_86 is signed(SUM_WIDTH_3_86-1 downto 0);
  constant SUM_WIDTH_3_87: positive := 9;
  subtype sum_t_3_87 is signed(SUM_WIDTH_3_87-1 downto 0);
  constant SUM_WIDTH_3_88: positive := 9;
  subtype sum_t_3_88 is signed(SUM_WIDTH_3_88-1 downto 0);
  constant SUM_WIDTH_3_89: positive := 9;
  subtype sum_t_3_89 is signed(SUM_WIDTH_3_89-1 downto 0);
  constant SUM_WIDTH_3_90: positive := 8;
  subtype sum_t_3_90 is signed(SUM_WIDTH_3_90-1 downto 0);
  constant SUM_WIDTH_3_91: positive := 9;
  subtype sum_t_3_91 is signed(SUM_WIDTH_3_91-1 downto 0);
  constant SUM_WIDTH_3_92: positive := 9;
  subtype sum_t_3_92 is signed(SUM_WIDTH_3_92-1 downto 0);
  constant SUM_WIDTH_3_93: positive := 9;
  subtype sum_t_3_93 is signed(SUM_WIDTH_3_93-1 downto 0);
  constant SUM_WIDTH_3_94: positive := 9;
  subtype sum_t_3_94 is signed(SUM_WIDTH_3_94-1 downto 0);
  constant SUM_WIDTH_3_95: positive := 9;
  subtype sum_t_3_95 is signed(SUM_WIDTH_3_95-1 downto 0);
  constant SUM_WIDTH_3_96: positive := 9;
  subtype sum_t_3_96 is signed(SUM_WIDTH_3_96-1 downto 0);
  constant SUM_WIDTH_3_97: positive := 8;
  subtype sum_t_3_97 is signed(SUM_WIDTH_3_97-1 downto 0);
  constant SUM_WIDTH_3_98: positive := 9;
  subtype sum_t_3_98 is signed(SUM_WIDTH_3_98-1 downto 0);
  constant SUM_WIDTH_3_99: positive := 7;
  subtype sum_t_3_99 is signed(SUM_WIDTH_3_99-1 downto 0);
  constant SUM_WIDTH_3_100: positive := 8;
  subtype sum_t_3_100 is signed(SUM_WIDTH_3_100-1 downto 0);
  constant SUM_WIDTH_3_101: positive := 9;
  subtype sum_t_3_101 is signed(SUM_WIDTH_3_101-1 downto 0);
  constant SUM_WIDTH_3_102: positive := 9;
  subtype sum_t_3_102 is signed(SUM_WIDTH_3_102-1 downto 0);
  constant SUM_WIDTH_3_103: positive := 9;
  subtype sum_t_3_103 is signed(SUM_WIDTH_3_103-1 downto 0);
  constant SUM_WIDTH_3_104: positive := 8;
  subtype sum_t_3_104 is signed(SUM_WIDTH_3_104-1 downto 0);
  constant SUM_WIDTH_3_105: positive := 8;
  subtype sum_t_3_105 is signed(SUM_WIDTH_3_105-1 downto 0);
  constant SUM_WIDTH_3_106: positive := 9;
  subtype sum_t_3_106 is signed(SUM_WIDTH_3_106-1 downto 0);
  constant SUM_WIDTH_3_107: positive := 9;
  subtype sum_t_3_107 is signed(SUM_WIDTH_3_107-1 downto 0);
  constant SUM_WIDTH_3_108: positive := 9;
  subtype sum_t_3_108 is signed(SUM_WIDTH_3_108-1 downto 0);
  constant SUM_WIDTH_3_109: positive := 9;
  subtype sum_t_3_109 is signed(SUM_WIDTH_3_109-1 downto 0);
  constant SUM_WIDTH_3_110: positive := 9;
  subtype sum_t_3_110 is signed(SUM_WIDTH_3_110-1 downto 0);
  constant SUM_WIDTH_3_111: positive := 8;
  subtype sum_t_3_111 is signed(SUM_WIDTH_3_111-1 downto 0);
  constant SUM_WIDTH_3_112: positive := 9;
  subtype sum_t_3_112 is signed(SUM_WIDTH_3_112-1 downto 0);
  constant SUM_WIDTH_3_113: positive := 9;
  subtype sum_t_3_113 is signed(SUM_WIDTH_3_113-1 downto 0);
  constant SUM_WIDTH_3_114: positive := 9;
  subtype sum_t_3_114 is signed(SUM_WIDTH_3_114-1 downto 0);
  constant SUM_WIDTH_3_115: positive := 9;
  subtype sum_t_3_115 is signed(SUM_WIDTH_3_115-1 downto 0);
  constant SUM_WIDTH_3_116: positive := 9;
  subtype sum_t_3_116 is signed(SUM_WIDTH_3_116-1 downto 0);
  constant SUM_WIDTH_3_117: positive := 8;
  subtype sum_t_3_117 is signed(SUM_WIDTH_3_117-1 downto 0);
  constant SUM_WIDTH_3_118: positive := 9;
  subtype sum_t_3_118 is signed(SUM_WIDTH_3_118-1 downto 0);
  constant SUM_WIDTH_3_119: positive := 9;
  subtype sum_t_3_119 is signed(SUM_WIDTH_3_119-1 downto 0);
  constant SUM_WIDTH_3_120: positive := 9;
  subtype sum_t_3_120 is signed(SUM_WIDTH_3_120-1 downto 0);
  constant SUM_WIDTH_3_121: positive := 8;
  subtype sum_t_3_121 is signed(SUM_WIDTH_3_121-1 downto 0);
  constant SUM_WIDTH_3_122: positive := 7;
  subtype sum_t_3_122 is signed(SUM_WIDTH_3_122-1 downto 0);
  constant SUM_WIDTH_3_123: positive := 9;
  subtype sum_t_3_123 is signed(SUM_WIDTH_3_123-1 downto 0);
  constant SUM_WIDTH_3_124: positive := 8;
  subtype sum_t_3_124 is signed(SUM_WIDTH_3_124-1 downto 0);
  constant SUM_WIDTH_3_125: positive := 8;
  subtype sum_t_3_125 is signed(SUM_WIDTH_3_125-1 downto 0);
  constant SUM_WIDTH_3_126: positive := 7;
  subtype sum_t_3_126 is signed(SUM_WIDTH_3_126-1 downto 0);
  constant SUM_WIDTH_3_127: positive := 8;
  subtype sum_t_3_127 is signed(SUM_WIDTH_3_127-1 downto 0);
  
  -- Function to saturate a signed value into W-bit signed range
  function saturate(x : signed; W : positive) return signed;
end package PkgKAN;

package body PkgKAN is
  -- Function to saturate a signed value into W-bit signed range
  function saturate(x : signed; W : positive) return signed is
      constant MAX_W_BITS : signed(W-1 downto 0) := (W-1 => '0', others => '1');
      constant MIN_W_BITS : signed(W-1 downto 0) := (W-1 => '1', others => '0');

      variable max_for_comp : signed(x'length-1 downto 0) := resize(MAX_W_BITS, x'length);
      variable min_for_comp : signed(x'length-1 downto 0) := resize(MIN_W_BITS, x'length);
      
      variable result : signed(W-1 downto 0);
  begin
      if x > max_for_comp then
          result := MAX_W_BITS;
      elsif x < min_for_comp then
          result := MIN_W_BITS;
      else
          result := resize(x, W);
      end if;

      return result;
  end function;
end package body PkgKAN;